magic
tech sky130A
magscale 1 2
timestamp 1608259780
<< metal1 >>
rect 8018 700612 8024 700664
rect 8076 700652 8082 700664
rect 8202 700652 8208 700664
rect 8076 700624 8208 700652
rect 8076 700612 8082 700624
rect 8202 700612 8208 700624
rect 8260 700652 8266 700664
rect 72970 700652 72976 700664
rect 8260 700624 72976 700652
rect 8260 700612 8266 700624
rect 72970 700612 72976 700624
rect 73028 700652 73034 700664
rect 137830 700652 137836 700664
rect 73028 700624 137836 700652
rect 73028 700612 73034 700624
rect 137830 700612 137836 700624
rect 137888 700652 137894 700664
rect 202782 700652 202788 700664
rect 137888 700624 202788 700652
rect 137888 700612 137894 700624
rect 202782 700612 202788 700624
rect 202840 700652 202846 700664
rect 267642 700652 267648 700664
rect 202840 700624 267648 700652
rect 202840 700612 202846 700624
rect 267642 700612 267648 700624
rect 267700 700612 267706 700664
rect 332502 700612 332508 700664
rect 332560 700652 332566 700664
rect 397454 700652 397460 700664
rect 332560 700624 397460 700652
rect 332560 700612 332566 700624
rect 397454 700612 397460 700624
rect 397512 700652 397518 700664
rect 462314 700652 462320 700664
rect 397512 700624 462320 700652
rect 397512 700612 397518 700624
rect 462314 700612 462320 700624
rect 462372 700652 462378 700664
rect 527174 700652 527180 700664
rect 462372 700624 527180 700652
rect 462372 700612 462378 700624
rect 527174 700612 527180 700624
rect 527232 700612 527238 700664
rect 272978 700272 272984 700324
rect 273036 700312 273042 700324
rect 283834 700312 283840 700324
rect 273036 700284 283840 700312
rect 273036 700272 273042 700284
rect 283834 700272 283840 700284
rect 283892 700272 283898 700324
rect 270862 700204 270868 700256
rect 270920 700244 270926 700256
rect 364978 700244 364984 700256
rect 270920 700216 364984 700244
rect 270920 700204 270926 700216
rect 364978 700204 364984 700216
rect 365036 700204 365042 700256
rect 218974 700136 218980 700188
rect 219032 700176 219038 700188
rect 312078 700176 312084 700188
rect 219032 700148 312084 700176
rect 219032 700136 219038 700148
rect 312078 700136 312084 700148
rect 312136 700136 312142 700188
rect 270678 700068 270684 700120
rect 270736 700108 270742 700120
rect 429838 700108 429844 700120
rect 270736 700080 429844 700108
rect 270736 700068 270742 700080
rect 429838 700068 429844 700080
rect 429896 700068 429902 700120
rect 89162 700000 89168 700052
rect 89220 700040 89226 700052
rect 312170 700040 312176 700052
rect 89220 700012 312176 700040
rect 89220 700000 89226 700012
rect 312170 700000 312176 700012
rect 312228 700000 312234 700052
rect 312722 700000 312728 700052
rect 312780 700040 312786 700052
rect 494790 700040 494796 700052
rect 312780 700012 494796 700040
rect 312780 700000 312786 700012
rect 494790 700000 494796 700012
rect 494848 700000 494854 700052
rect 154114 699932 154120 699984
rect 154172 699972 154178 699984
rect 268562 699972 268568 699984
rect 154172 699944 268568 699972
rect 154172 699932 154178 699944
rect 268562 699932 268568 699944
rect 268620 699932 268626 699984
rect 270770 699932 270776 699984
rect 270828 699972 270834 699984
rect 559650 699972 559656 699984
rect 270828 699944 559656 699972
rect 270828 699932 270834 699944
rect 559650 699932 559656 699944
rect 559708 699932 559714 699984
rect 24302 699864 24308 699916
rect 24360 699904 24366 699916
rect 314470 699904 314476 699916
rect 24360 699876 314476 699904
rect 24360 699864 24366 699876
rect 314470 699864 314476 699876
rect 314528 699864 314534 699916
rect 527174 699864 527180 699916
rect 527232 699904 527238 699916
rect 579890 699904 579896 699916
rect 527232 699876 579896 699904
rect 527232 699864 527238 699876
rect 579890 699864 579896 699876
rect 579948 699864 579954 699916
rect 561490 674160 561496 674212
rect 561548 674200 561554 674212
rect 578510 674200 578516 674212
rect 561548 674172 578516 674200
rect 561548 674160 561554 674172
rect 578510 674160 578516 674172
rect 578568 674160 578574 674212
rect 2958 653488 2964 653540
rect 3016 653528 3022 653540
rect 8018 653528 8024 653540
rect 3016 653500 8024 653528
rect 3016 653488 3022 653500
rect 8018 653488 8024 653500
rect 8076 653488 8082 653540
rect 270494 627104 270500 627156
rect 270552 627144 270558 627156
rect 578786 627144 578792 627156
rect 270552 627116 578792 627144
rect 270552 627104 270558 627116
rect 578786 627104 578792 627116
rect 578844 627104 578850 627156
rect 49602 586576 49608 586628
rect 49660 586616 49666 586628
rect 313734 586616 313740 586628
rect 49660 586588 313740 586616
rect 49660 586576 49666 586588
rect 313734 586576 313740 586588
rect 313792 586576 313798 586628
rect 217962 586508 217968 586560
rect 218020 586548 218026 586560
rect 270586 586548 270592 586560
rect 218020 586520 270592 586548
rect 218020 586508 218026 586520
rect 270586 586508 270592 586520
rect 270644 586548 270650 586560
rect 271138 586548 271144 586560
rect 270644 586520 271144 586548
rect 270644 586508 270650 586520
rect 271138 586508 271144 586520
rect 271196 586508 271202 586560
rect 306190 586508 306196 586560
rect 306248 586548 306254 586560
rect 316402 586548 316408 586560
rect 306248 586520 316408 586548
rect 306248 586508 306254 586520
rect 316402 586508 316408 586520
rect 316460 586508 316466 586560
rect 326890 586508 326896 586560
rect 326948 586548 326954 586560
rect 337010 586548 337016 586560
rect 326948 586520 337016 586548
rect 326948 586508 326954 586520
rect 337010 586508 337016 586520
rect 337068 586508 337074 586560
rect 347406 586508 347412 586560
rect 347464 586548 347470 586560
rect 357618 586548 357624 586560
rect 347464 586520 357624 586548
rect 347464 586508 347470 586520
rect 357618 586508 357624 586520
rect 357676 586508 357682 586560
rect 73522 586440 73528 586492
rect 73580 586480 73586 586492
rect 272242 586480 272248 586492
rect 73580 586452 272248 586480
rect 73580 586440 73586 586452
rect 272242 586440 272248 586452
rect 272300 586480 272306 586492
rect 365438 586480 365444 586492
rect 272300 586452 365444 586480
rect 272300 586440 272306 586452
rect 365438 586440 365444 586452
rect 365496 586440 365502 586492
rect 368014 586440 368020 586492
rect 368072 586480 368078 586492
rect 378226 586480 378232 586492
rect 368072 586452 378232 586480
rect 368072 586440 368078 586452
rect 378226 586440 378232 586452
rect 378284 586440 378290 586492
rect 388622 586440 388628 586492
rect 388680 586480 388686 586492
rect 398834 586480 398840 586492
rect 388680 586452 398840 586480
rect 388680 586440 388686 586452
rect 398834 586440 398840 586452
rect 398892 586440 398898 586492
rect 409230 586440 409236 586492
rect 409288 586480 409294 586492
rect 415118 586480 415124 586492
rect 409288 586452 415124 586480
rect 409288 586440 409294 586452
rect 415118 586440 415124 586452
rect 415176 586440 415182 586492
rect 463694 586480 463700 586492
rect 458468 586452 463700 586480
rect 242066 586372 242072 586424
rect 242124 586412 242130 586424
rect 292942 586412 292948 586424
rect 242124 586384 292948 586412
rect 242124 586372 242130 586384
rect 292942 586372 292948 586384
rect 293000 586372 293006 586424
rect 300210 586372 300216 586424
rect 300268 586412 300274 586424
rect 437750 586412 437756 586424
rect 300268 586384 437756 586412
rect 300268 586372 300274 586384
rect 437750 586372 437756 586384
rect 437808 586372 437814 586424
rect 456242 586412 456248 586424
rect 445956 586384 456248 586412
rect 169754 586304 169760 586356
rect 169812 586344 169818 586356
rect 313642 586344 313648 586356
rect 169812 586316 313648 586344
rect 169812 586304 169818 586316
rect 313642 586304 313648 586316
rect 313700 586304 313706 586356
rect 313734 586304 313740 586356
rect 313792 586344 313798 586356
rect 341518 586344 341524 586356
rect 313792 586316 341524 586344
rect 313792 586304 313798 586316
rect 341518 586304 341524 586316
rect 341576 586304 341582 586356
rect 121730 586236 121736 586288
rect 121788 586276 121794 586288
rect 312354 586276 312360 586288
rect 121788 586248 312360 586276
rect 121788 586236 121794 586248
rect 312354 586236 312360 586248
rect 312412 586236 312418 586288
rect 312814 586236 312820 586288
rect 312872 586276 312878 586288
rect 413646 586276 413652 586288
rect 312872 586248 413652 586276
rect 312872 586236 312878 586248
rect 413646 586236 413652 586248
rect 413704 586236 413710 586288
rect 415118 586236 415124 586288
rect 415176 586276 415182 586288
rect 415176 586248 425376 586276
rect 415176 586236 415182 586248
rect 198734 586168 198740 586220
rect 198792 586208 198798 586220
rect 209038 586208 209044 586220
rect 198792 586180 209044 586208
rect 198792 586168 198798 586180
rect 209038 586168 209044 586180
rect 209096 586168 209102 586220
rect 216490 586168 216496 586220
rect 216548 586208 216554 586220
rect 229646 586208 229652 586220
rect 216548 586180 229652 586208
rect 216548 586168 216554 586180
rect 229646 586168 229652 586180
rect 229704 586168 229710 586220
rect 306190 586208 306196 586220
rect 270512 586180 306196 586208
rect 239950 586100 239956 586152
rect 240008 586140 240014 586152
rect 250254 586140 250260 586152
rect 240008 586112 250260 586140
rect 240008 586100 240014 586112
rect 250254 586100 250260 586112
rect 250312 586100 250318 586152
rect 270402 586140 270408 586152
rect 267936 586112 270408 586140
rect 145834 586032 145840 586084
rect 145892 586072 145898 586084
rect 267090 586072 267096 586084
rect 145892 586044 267096 586072
rect 145892 586032 145898 586044
rect 267090 586032 267096 586044
rect 267148 586032 267154 586084
rect 193858 585964 193864 586016
rect 193916 586004 193922 586016
rect 198734 586004 198740 586016
rect 193916 585976 198740 586004
rect 193916 585964 193922 585976
rect 198734 585964 198740 585976
rect 198792 585964 198798 586016
rect 229646 585964 229652 586016
rect 229704 586004 229710 586016
rect 229704 585976 239904 586004
rect 229704 585964 229710 585976
rect 209038 585896 209044 585948
rect 209096 585936 209102 585948
rect 216398 585936 216404 585948
rect 209096 585908 216404 585936
rect 209096 585896 209102 585908
rect 216398 585896 216404 585908
rect 216456 585896 216462 585948
rect 239876 585936 239904 585976
rect 257614 585964 257620 586016
rect 257672 585964 257678 586016
rect 267734 585964 267740 586016
rect 267792 586004 267798 586016
rect 267936 586004 267964 586112
rect 270402 586100 270408 586112
rect 270460 586140 270466 586152
rect 270512 586140 270540 586180
rect 306190 586168 306196 586180
rect 306248 586168 306254 586220
rect 316402 586168 316408 586220
rect 316460 586208 316466 586220
rect 326890 586208 326896 586220
rect 316460 586180 326896 586208
rect 316460 586168 316466 586180
rect 326890 586168 326896 586180
rect 326948 586168 326954 586220
rect 337010 586168 337016 586220
rect 337068 586208 337074 586220
rect 347406 586208 347412 586220
rect 337068 586180 347412 586208
rect 337068 586168 337074 586180
rect 347406 586168 347412 586180
rect 347464 586168 347470 586220
rect 357618 586168 357624 586220
rect 357676 586208 357682 586220
rect 368014 586208 368020 586220
rect 357676 586180 368020 586208
rect 357676 586168 357682 586180
rect 368014 586168 368020 586180
rect 368072 586168 368078 586220
rect 378226 586168 378232 586220
rect 378284 586208 378290 586220
rect 388622 586208 388628 586220
rect 378284 586180 388628 586208
rect 378284 586168 378290 586180
rect 388622 586168 388628 586180
rect 388680 586168 388686 586220
rect 398834 586168 398840 586220
rect 398892 586208 398898 586220
rect 409230 586208 409236 586220
rect 398892 586180 409236 586208
rect 398892 586168 398898 586180
rect 409230 586168 409236 586180
rect 409288 586168 409294 586220
rect 425348 586208 425376 586248
rect 442994 586236 443000 586288
rect 443052 586276 443058 586288
rect 445956 586276 445984 586384
rect 456242 586372 456248 586384
rect 456300 586372 456306 586424
rect 456334 586372 456340 586424
rect 456392 586412 456398 586424
rect 458468 586412 458496 586452
rect 463694 586440 463700 586452
rect 463752 586440 463758 586492
rect 485774 586480 485780 586492
rect 479076 586452 485780 586480
rect 456392 586384 458496 586412
rect 456392 586372 456398 586384
rect 473906 586372 473912 586424
rect 473964 586412 473970 586424
rect 476850 586412 476856 586424
rect 473964 586384 476856 586412
rect 473964 586372 473970 586384
rect 476850 586372 476856 586384
rect 476908 586372 476914 586424
rect 476942 586372 476948 586424
rect 477000 586412 477006 586424
rect 479076 586412 479104 586452
rect 485774 586440 485780 586452
rect 485832 586440 485838 586492
rect 477000 586384 479104 586412
rect 477000 586372 477006 586384
rect 443052 586248 445984 586276
rect 443052 586236 443058 586248
rect 432782 586208 432788 586220
rect 425348 586180 432788 586208
rect 432782 586168 432788 586180
rect 432840 586168 432846 586220
rect 270460 586112 270540 586140
rect 270460 586100 270466 586112
rect 292942 586100 292948 586152
rect 293000 586140 293006 586152
rect 294322 586140 294328 586152
rect 293000 586112 294328 586140
rect 293000 586100 293006 586112
rect 294322 586100 294328 586112
rect 294380 586140 294386 586152
rect 533982 586140 533988 586152
rect 294380 586112 533988 586140
rect 294380 586100 294386 586112
rect 533982 586100 533988 586112
rect 534040 586100 534046 586152
rect 271138 586032 271144 586084
rect 271196 586072 271202 586084
rect 509878 586072 509884 586084
rect 271196 586044 509884 586072
rect 271196 586032 271202 586044
rect 509878 586032 509884 586044
rect 509936 586032 509942 586084
rect 267792 585976 267964 586004
rect 270328 585976 270540 586004
rect 267792 585964 267798 585976
rect 239950 585936 239956 585948
rect 239876 585908 239956 585936
rect 239950 585896 239956 585908
rect 240008 585896 240014 585948
rect 250254 585896 250260 585948
rect 250312 585936 250318 585948
rect 257632 585936 257660 585964
rect 250312 585908 257660 585936
rect 250312 585896 250318 585908
rect 265986 585896 265992 585948
rect 266044 585936 266050 585948
rect 270328 585936 270356 585976
rect 266044 585908 270356 585936
rect 270512 585936 270540 585976
rect 313642 585964 313648 586016
rect 313700 586004 313706 586016
rect 461670 586004 461676 586016
rect 313700 585976 461676 586004
rect 313700 585964 313706 585976
rect 461670 585964 461676 585976
rect 461728 585964 461734 586016
rect 288526 585936 288532 585948
rect 270512 585908 288532 585936
rect 266044 585896 266050 585908
rect 288526 585896 288532 585908
rect 288584 585936 288590 585948
rect 557902 585936 557908 585948
rect 288584 585908 557908 585936
rect 288584 585896 288590 585908
rect 557902 585896 557908 585908
rect 557960 585896 557966 585948
rect 318610 582904 318616 582956
rect 318668 582944 318674 582956
rect 560846 582944 560852 582956
rect 318668 582916 560852 582944
rect 318668 582904 318674 582916
rect 560846 582904 560852 582916
rect 560904 582904 560910 582956
rect 26510 582360 26516 582412
rect 26568 582400 26574 582412
rect 270034 582400 270040 582412
rect 26568 582372 270040 582400
rect 26568 582360 26574 582372
rect 270034 582360 270040 582372
rect 270092 582360 270098 582412
rect 27246 582292 27252 582344
rect 27304 582332 27310 582344
rect 275922 582332 275928 582344
rect 27304 582304 275928 582332
rect 27304 582292 27310 582304
rect 275922 582292 275928 582304
rect 275980 582292 275986 582344
rect 24854 582224 24860 582276
rect 24912 582264 24918 582276
rect 314286 582264 314292 582276
rect 24912 582236 314292 582264
rect 24912 582224 24918 582236
rect 314286 582224 314292 582236
rect 314344 582224 314350 582276
rect 319438 582224 319444 582276
rect 319496 582264 319502 582276
rect 558454 582264 558460 582276
rect 319496 582236 558460 582264
rect 319496 582224 319502 582236
rect 558454 582224 558460 582236
rect 558512 582224 558518 582276
rect 275922 580660 275928 580712
rect 275980 580700 275986 580712
rect 315022 580700 315028 580712
rect 275980 580672 315028 580700
rect 275980 580660 275986 580672
rect 315022 580660 315028 580672
rect 315080 580660 315086 580712
rect 26510 577096 26516 577108
rect 25056 577068 26516 577096
rect 24946 576988 24952 577040
rect 25004 577028 25010 577040
rect 25056 577028 25084 577068
rect 26510 577056 26516 577068
rect 26568 577056 26574 577108
rect 25004 577000 25084 577028
rect 25004 576988 25010 577000
rect 317966 576240 317972 576292
rect 318024 576280 318030 576292
rect 319438 576280 319444 576292
rect 318024 576252 319444 576280
rect 318024 576240 318030 576252
rect 319438 576240 319444 576252
rect 319496 576240 319502 576292
rect 317138 572636 317144 572688
rect 317196 572676 317202 572688
rect 317966 572676 317972 572688
rect 317196 572648 317972 572676
rect 317196 572636 317202 572648
rect 317966 572636 317972 572648
rect 318024 572636 318030 572688
rect 270034 569576 270040 569628
rect 270092 569616 270098 569628
rect 273806 569616 273812 569628
rect 270092 569588 273812 569616
rect 270092 569576 270098 569588
rect 273806 569576 273812 569588
rect 273864 569576 273870 569628
rect 273806 565836 273812 565888
rect 273864 565876 273870 565888
rect 275278 565876 275284 565888
rect 273864 565848 275284 565876
rect 273864 565836 273870 565848
rect 275278 565836 275284 565848
rect 275336 565836 275342 565888
rect 275278 562776 275284 562828
rect 275336 562816 275342 562828
rect 279602 562816 279608 562828
rect 275336 562788 279608 562816
rect 275336 562776 275342 562788
rect 279602 562776 279608 562788
rect 279660 562776 279666 562828
rect 315022 562300 315028 562352
rect 315080 562340 315086 562352
rect 317138 562340 317144 562352
rect 315080 562312 317144 562340
rect 315080 562300 315086 562312
rect 317138 562300 317144 562312
rect 317196 562300 317202 562352
rect 315022 559416 315028 559428
rect 312096 559388 315028 559416
rect 309778 559308 309784 559360
rect 309836 559348 309842 559360
rect 312096 559348 312124 559388
rect 315022 559376 315028 559388
rect 315080 559376 315086 559428
rect 309836 559320 312124 559348
rect 309836 559308 309842 559320
rect 279694 556452 279700 556504
rect 279752 556492 279758 556504
rect 279752 556464 282684 556492
rect 279752 556452 279758 556464
rect 282656 556424 282684 556464
rect 285490 556424 285496 556436
rect 282656 556396 285496 556424
rect 285490 556384 285496 556396
rect 285548 556384 285554 556436
rect 285490 549720 285496 549772
rect 285548 549760 285554 549772
rect 290642 549760 290648 549772
rect 285548 549732 290648 549760
rect 285548 549720 285554 549732
rect 290642 549720 290648 549732
rect 290700 549720 290706 549772
rect 269298 547612 269304 547664
rect 269356 547652 269362 547664
rect 269356 547624 313596 547652
rect 269356 547612 269362 547624
rect 313568 547584 313596 547624
rect 314194 547584 314200 547596
rect 313568 547556 314200 547584
rect 314194 547544 314200 547556
rect 314252 547584 314258 547596
rect 318610 547584 318616 547596
rect 314252 547556 318616 547584
rect 314252 547544 314258 547556
rect 318610 547544 318616 547556
rect 318668 547544 318674 547596
rect 314286 544892 314292 544944
rect 314344 544932 314350 544944
rect 315022 544932 315028 544944
rect 314344 544904 315028 544932
rect 314344 544892 314350 544904
rect 315022 544892 315028 544904
rect 315080 544892 315086 544944
rect 307662 544552 307668 544604
rect 307720 544592 307726 544604
rect 309778 544592 309784 544604
rect 307720 544564 309784 544592
rect 307720 544552 307726 544564
rect 309778 544552 309784 544564
rect 309836 544552 309842 544604
rect 290642 540200 290648 540252
rect 290700 540240 290706 540252
rect 290700 540212 291516 540240
rect 290700 540200 290706 540212
rect 291488 540172 291516 540212
rect 293310 540172 293316 540184
rect 291488 540144 293316 540172
rect 293310 540132 293316 540144
rect 293368 540132 293374 540184
rect 293310 537208 293316 537260
rect 293368 537248 293374 537260
rect 294414 537248 294420 537260
rect 293368 537220 294420 537248
rect 293368 537208 293374 537220
rect 294414 537208 294420 537220
rect 294472 537208 294478 537260
rect 304718 536528 304724 536580
rect 304776 536568 304782 536580
rect 307662 536568 307668 536580
rect 304776 536540 307668 536568
rect 304776 536528 304782 536540
rect 307662 536528 307668 536540
rect 307720 536528 307726 536580
rect 303246 534488 303252 534540
rect 303304 534528 303310 534540
rect 304718 534528 304724 534540
rect 303304 534500 304724 534528
rect 303304 534488 303310 534500
rect 304718 534488 304724 534500
rect 304776 534488 304782 534540
rect 294414 534352 294420 534404
rect 294472 534392 294478 534404
rect 294472 534364 295932 534392
rect 294472 534352 294478 534364
rect 295904 534256 295932 534364
rect 298002 534256 298008 534268
rect 295904 534228 298008 534256
rect 298002 534216 298008 534228
rect 298060 534216 298066 534268
rect 303246 529972 303252 529984
rect 300320 529944 303252 529972
rect 298830 529864 298836 529916
rect 298888 529904 298894 529916
rect 300320 529904 300348 529944
rect 303246 529932 303252 529944
rect 303304 529932 303310 529984
rect 298888 529876 300348 529904
rect 298888 529864 298894 529876
rect 298002 523948 298008 524000
rect 298060 523988 298066 524000
rect 300118 523988 300124 524000
rect 298060 523960 300124 523988
rect 298060 523948 298066 523960
rect 300118 523948 300124 523960
rect 300176 523948 300182 524000
rect 295058 522588 295064 522640
rect 295116 522628 295122 522640
rect 298738 522628 298744 522640
rect 295116 522600 298744 522628
rect 295116 522588 295122 522600
rect 298738 522588 298744 522600
rect 298796 522588 298802 522640
rect 300118 519052 300124 519104
rect 300176 519092 300182 519104
rect 301590 519092 301596 519104
rect 300176 519064 301596 519092
rect 300176 519052 300182 519064
rect 301590 519052 301596 519064
rect 301648 519052 301654 519104
rect 301590 516672 301596 516724
rect 301648 516712 301654 516724
rect 303154 516712 303160 516724
rect 301648 516684 303160 516712
rect 301648 516672 301654 516684
rect 303154 516672 303160 516684
rect 303212 516672 303218 516724
rect 303154 515176 303160 515228
rect 303212 515216 303218 515228
rect 303212 515188 306144 515216
rect 303212 515176 303218 515188
rect 306116 515148 306144 515188
rect 307386 515148 307392 515160
rect 306116 515120 307392 515148
rect 307386 515108 307392 515120
rect 307444 515108 307450 515160
rect 558454 512116 558460 512168
rect 558512 512156 558518 512168
rect 558914 512156 558920 512168
rect 558512 512128 558920 512156
rect 558512 512116 558518 512128
rect 558914 512116 558920 512128
rect 558972 512116 558978 512168
rect 269298 511504 269304 511556
rect 269356 511544 269362 511556
rect 272150 511544 272156 511556
rect 269356 511516 272156 511544
rect 269356 511504 269362 511516
rect 272150 511504 272156 511516
rect 272208 511544 272214 511556
rect 295058 511544 295064 511556
rect 272208 511516 295064 511544
rect 272208 511504 272214 511516
rect 295058 511504 295064 511516
rect 295116 511504 295122 511556
rect 307386 509668 307392 509720
rect 307444 509708 307450 509720
rect 315022 509708 315028 509720
rect 307444 509680 315028 509708
rect 307444 509668 307450 509680
rect 315022 509668 315028 509680
rect 315080 509668 315086 509720
rect 307386 487228 307392 487280
rect 307444 487268 307450 487280
rect 307570 487268 307576 487280
rect 307444 487240 307576 487268
rect 307444 487228 307450 487240
rect 307570 487228 307576 487240
rect 307628 487228 307634 487280
rect 2958 479884 2964 479936
rect 3016 479924 3022 479936
rect 3970 479924 3976 479936
rect 3016 479896 3976 479924
rect 3016 479884 3022 479896
rect 3970 479884 3976 479896
rect 4028 479884 4034 479936
rect 270034 472540 270040 472592
rect 270092 472580 270098 472592
rect 315022 472580 315028 472592
rect 270092 472552 315028 472580
rect 270092 472540 270098 472552
rect 315022 472540 315028 472552
rect 315080 472540 315086 472592
rect 307386 466624 307392 466676
rect 307444 466664 307450 466676
rect 307570 466664 307576 466676
rect 307444 466636 307576 466664
rect 307444 466624 307450 466636
rect 307570 466624 307576 466636
rect 307628 466624 307634 466676
rect 307386 446020 307392 446072
rect 307444 446060 307450 446072
rect 307570 446060 307576 446072
rect 307444 446032 307576 446060
rect 307444 446020 307450 446032
rect 307570 446020 307576 446032
rect 307628 446020 307634 446072
rect 558454 440444 558460 440496
rect 558512 440484 558518 440496
rect 558914 440484 558920 440496
rect 558512 440456 558920 440484
rect 558512 440444 558518 440456
rect 558914 440444 558920 440456
rect 558972 440444 558978 440496
rect 269298 440104 269304 440156
rect 269356 440144 269362 440156
rect 286226 440144 286232 440156
rect 269356 440116 286232 440144
rect 269356 440104 269362 440116
rect 286226 440104 286232 440116
rect 286284 440104 286290 440156
rect 307386 425416 307392 425468
rect 307444 425456 307450 425468
rect 307570 425456 307576 425468
rect 307444 425428 307576 425456
rect 307444 425416 307450 425428
rect 307570 425416 307576 425428
rect 307628 425416 307634 425468
rect 269298 404812 269304 404864
rect 269356 404852 269362 404864
rect 303890 404852 303896 404864
rect 269356 404824 303896 404852
rect 269356 404812 269362 404824
rect 303890 404812 303896 404824
rect 303948 404812 303954 404864
rect 298756 386464 298876 386492
rect 298756 386436 298784 386464
rect 298848 386436 298876 386464
rect 298738 386384 298744 386436
rect 298796 386384 298802 386436
rect 298830 386384 298836 386436
rect 298888 386384 298894 386436
rect 291378 386356 291384 386368
rect 41156 386328 44036 386356
rect 24946 386180 24952 386232
rect 25004 386220 25010 386232
rect 41156 386220 41184 386328
rect 25004 386192 30972 386220
rect 25004 386180 25010 386192
rect 30944 385948 30972 386192
rect 33888 386192 41184 386220
rect 44008 386220 44036 386328
rect 56612 386328 61976 386356
rect 56612 386220 56640 386328
rect 44008 386192 56640 386220
rect 61948 386220 61976 386328
rect 77220 386328 82584 386356
rect 77220 386220 77248 386328
rect 61948 386192 77248 386220
rect 82556 386220 82584 386328
rect 97828 386328 103284 386356
rect 97828 386220 97856 386328
rect 82556 386192 97856 386220
rect 103256 386220 103284 386328
rect 123588 386328 126468 386356
rect 123588 386220 123616 386328
rect 103256 386192 113404 386220
rect 33888 385948 33916 386192
rect 30944 385920 33916 385948
rect 113376 385948 113404 386192
rect 116320 386192 123616 386220
rect 126440 386220 126468 386328
rect 144196 386328 147076 386356
rect 144196 386220 144224 386328
rect 126440 386192 134012 386220
rect 116320 385948 116348 386192
rect 113376 385920 116348 385948
rect 133984 385948 134012 386192
rect 136928 386192 144224 386220
rect 147048 386220 147076 386328
rect 164804 386328 167868 386356
rect 164804 386220 164832 386328
rect 167840 386288 167868 386328
rect 190564 386328 198596 386356
rect 167840 386260 178080 386288
rect 147048 386192 154620 386220
rect 136928 385948 136956 386192
rect 133984 385920 136956 385948
rect 154592 385948 154620 386192
rect 157536 386192 164832 386220
rect 178052 386220 178080 386260
rect 190564 386220 190592 386328
rect 198568 386288 198596 386328
rect 247236 386328 250300 386356
rect 198568 386260 211200 386288
rect 178052 386192 190592 386220
rect 211172 386220 211200 386260
rect 226628 386260 231854 386288
rect 226628 386220 226656 386260
rect 211172 386192 216444 386220
rect 157536 385948 157564 386192
rect 154592 385920 157564 385948
rect 216416 385948 216444 386192
rect 219360 386192 226656 386220
rect 231826 386220 231854 386260
rect 247236 386220 247264 386328
rect 250272 386288 250300 386328
rect 281092 386328 291384 386356
rect 250272 386260 260512 386288
rect 231826 386192 237052 386220
rect 219360 385948 219388 386192
rect 216416 385920 219388 385948
rect 237024 385948 237052 386192
rect 239968 386192 247264 386220
rect 260484 386220 260512 386260
rect 278130 386248 278136 386300
rect 278188 386288 278194 386300
rect 281092 386288 281120 386328
rect 291378 386316 291384 386328
rect 291436 386316 291442 386368
rect 309042 386316 309048 386368
rect 309100 386356 309106 386368
rect 314378 386356 314384 386368
rect 309100 386328 314384 386356
rect 309100 386316 309106 386328
rect 314378 386316 314384 386328
rect 314436 386316 314442 386368
rect 278188 386260 281120 386288
rect 278188 386248 278194 386260
rect 286226 386248 286232 386300
rect 286284 386288 286290 386300
rect 558454 386288 558460 386300
rect 286284 386260 558460 386288
rect 286284 386248 286290 386260
rect 558454 386248 558460 386260
rect 558512 386248 558518 386300
rect 267918 386220 267924 386232
rect 260484 386192 267924 386220
rect 239968 385948 239996 386192
rect 267918 386180 267924 386192
rect 267976 386180 267982 386232
rect 291378 386112 291384 386164
rect 291436 386152 291442 386164
rect 298738 386152 298744 386164
rect 291436 386124 298744 386152
rect 291436 386112 291442 386124
rect 298738 386112 298744 386124
rect 298796 386112 298802 386164
rect 237024 385920 239996 385948
rect 314010 385704 314016 385756
rect 314068 385744 314074 385756
rect 314378 385744 314384 385756
rect 314068 385716 314384 385744
rect 314068 385704 314074 385716
rect 314378 385704 314384 385716
rect 314436 385704 314442 385756
rect 303890 384888 303896 384940
rect 303948 384928 303954 384940
rect 312630 384928 312636 384940
rect 303948 384900 312636 384928
rect 303948 384888 303954 384900
rect 312630 384888 312636 384900
rect 312688 384928 312694 384940
rect 560846 384928 560852 384940
rect 312688 384900 560852 384928
rect 312688 384888 312694 384900
rect 560846 384888 560852 384900
rect 560904 384888 560910 384940
rect 307386 384208 307392 384260
rect 307444 384248 307450 384260
rect 307570 384248 307576 384260
rect 307444 384220 307576 384248
rect 307444 384208 307450 384220
rect 307570 384208 307576 384220
rect 307628 384208 307634 384260
rect 256050 382644 256056 382696
rect 256108 382684 256114 382696
rect 271046 382684 271052 382696
rect 256108 382656 271052 382684
rect 256108 382644 256114 382656
rect 271046 382644 271052 382656
rect 271104 382644 271110 382696
rect 275278 382644 275284 382696
rect 275336 382684 275342 382696
rect 286318 382684 286324 382696
rect 275336 382656 286324 382684
rect 275336 382644 275342 382656
rect 286318 382644 286324 382656
rect 286376 382644 286382 382696
rect 301682 382644 301688 382696
rect 301740 382684 301746 382696
rect 331490 382684 331496 382696
rect 301740 382656 331496 382684
rect 301740 382644 301746 382656
rect 331490 382644 331496 382656
rect 331548 382644 331554 382696
rect 232130 382576 232136 382628
rect 232188 382616 232194 382628
rect 313550 382616 313556 382628
rect 232188 382588 313556 382616
rect 232188 382576 232194 382588
rect 313550 382576 313556 382588
rect 313608 382576 313614 382628
rect 270126 382508 270132 382560
rect 270184 382548 270190 382560
rect 355594 382548 355600 382560
rect 270184 382520 355600 382548
rect 270184 382508 270190 382520
rect 355594 382508 355600 382520
rect 355652 382508 355658 382560
rect 270954 382440 270960 382492
rect 271012 382480 271018 382492
rect 271966 382480 271972 382492
rect 271012 382452 271972 382480
rect 271012 382440 271018 382452
rect 271966 382440 271972 382452
rect 272024 382480 272030 382492
rect 379514 382480 379520 382492
rect 272024 382452 379520 382480
rect 272024 382440 272030 382452
rect 379514 382440 379520 382452
rect 379572 382440 379578 382492
rect 208026 382372 208032 382424
rect 208084 382412 208090 382424
rect 278222 382412 278228 382424
rect 208084 382384 278228 382412
rect 208084 382372 208090 382384
rect 278222 382372 278228 382384
rect 278280 382412 278286 382424
rect 279510 382412 279516 382424
rect 278280 382384 279516 382412
rect 278280 382372 278286 382384
rect 279510 382372 279516 382384
rect 279568 382372 279574 382424
rect 279694 382372 279700 382424
rect 279752 382412 279758 382424
rect 403618 382412 403624 382424
rect 279752 382384 403624 382412
rect 279752 382372 279758 382384
rect 403618 382372 403624 382384
rect 403676 382372 403682 382424
rect 183922 382304 183928 382356
rect 183980 382344 183986 382356
rect 264974 382344 264980 382356
rect 183980 382316 264980 382344
rect 183980 382304 183986 382316
rect 264974 382304 264980 382316
rect 265032 382304 265038 382356
rect 275186 382304 275192 382356
rect 275244 382344 275250 382356
rect 275278 382344 275284 382356
rect 275244 382316 275284 382344
rect 275244 382304 275250 382316
rect 275278 382304 275284 382316
rect 275336 382304 275342 382356
rect 111794 382236 111800 382288
rect 111852 382276 111858 382288
rect 279694 382276 279700 382288
rect 111852 382248 279700 382276
rect 111852 382236 111858 382248
rect 279694 382236 279700 382248
rect 279752 382236 279758 382288
rect 286318 382236 286324 382288
rect 286376 382276 286382 382288
rect 295886 382276 295892 382288
rect 286376 382248 295892 382276
rect 286376 382236 286382 382248
rect 295886 382236 295892 382248
rect 295944 382236 295950 382288
rect 316402 382236 316408 382288
rect 316460 382276 316466 382288
rect 475930 382276 475936 382288
rect 316460 382248 475936 382276
rect 316460 382236 316466 382248
rect 475930 382236 475936 382248
rect 475988 382236 475994 382288
rect 135898 382168 135904 382220
rect 135956 382208 135962 382220
rect 314102 382208 314108 382220
rect 135956 382180 314108 382208
rect 135956 382168 135962 382180
rect 314102 382168 314108 382180
rect 314160 382208 314166 382220
rect 427722 382208 427728 382220
rect 314160 382180 427728 382208
rect 314160 382168 314166 382180
rect 427722 382168 427728 382180
rect 427780 382168 427786 382220
rect 87690 382100 87696 382152
rect 87748 382140 87754 382152
rect 270954 382140 270960 382152
rect 87748 382112 270960 382140
rect 87748 382100 87754 382112
rect 270954 382100 270960 382112
rect 271012 382100 271018 382152
rect 279510 382100 279516 382152
rect 279568 382140 279574 382152
rect 499850 382140 499856 382152
rect 279568 382112 499856 382140
rect 279568 382100 279574 382112
rect 499850 382100 499856 382112
rect 499908 382100 499914 382152
rect 39666 382032 39672 382084
rect 39724 382072 39730 382084
rect 301682 382072 301688 382084
rect 39724 382044 301688 382072
rect 39724 382032 39730 382044
rect 301682 382032 301688 382044
rect 301740 382032 301746 382084
rect 313550 382032 313556 382084
rect 313608 382072 313614 382084
rect 313918 382072 313924 382084
rect 313608 382044 313924 382072
rect 313608 382032 313614 382044
rect 313918 382032 313924 382044
rect 313976 382072 313982 382084
rect 523954 382072 523960 382084
rect 313976 382044 523960 382072
rect 313976 382032 313982 382044
rect 523954 382032 523960 382044
rect 524012 382032 524018 382084
rect 63770 381964 63776 382016
rect 63828 382004 63834 382016
rect 270126 382004 270132 382016
rect 63828 381976 270132 382004
rect 63828 381964 63834 381976
rect 270126 381964 270132 381976
rect 270184 381964 270190 382016
rect 271046 381964 271052 382016
rect 271104 382004 271110 382016
rect 272058 382004 272064 382016
rect 271104 381976 272064 382004
rect 271104 381964 271110 381976
rect 272058 381964 272064 381976
rect 272116 382004 272122 382016
rect 548058 382004 548064 382016
rect 272116 381976 548064 382004
rect 272116 381964 272122 381976
rect 548058 381964 548064 381976
rect 548116 381964 548122 382016
rect 264974 381896 264980 381948
rect 265032 381936 265038 381948
rect 275186 381936 275192 381948
rect 265032 381908 275192 381936
rect 265032 381896 265038 381908
rect 275186 381896 275192 381908
rect 275244 381896 275250 381948
rect 295886 381896 295892 381948
rect 295944 381936 295950 381948
rect 313826 381936 313832 381948
rect 295944 381908 313832 381936
rect 295944 381896 295950 381908
rect 313826 381896 313832 381908
rect 313884 381936 313890 381948
rect 316402 381936 316408 381948
rect 313884 381908 316408 381936
rect 313884 381896 313890 381908
rect 316402 381896 316408 381908
rect 316460 381896 316466 381948
rect 273162 359388 273168 359440
rect 273220 359428 273226 359440
rect 278590 359428 278596 359440
rect 273220 359400 278596 359428
rect 273220 359388 273226 359400
rect 278590 359388 278596 359400
rect 278648 359388 278654 359440
rect 306926 359428 306932 359440
rect 301792 359400 306932 359428
rect 273346 359320 273352 359372
rect 273404 359360 273410 359372
rect 286226 359360 286232 359372
rect 273404 359332 286232 359360
rect 273404 359320 273410 359332
rect 286226 359320 286232 359332
rect 286284 359320 286290 359372
rect 301222 359320 301228 359372
rect 301280 359360 301286 359372
rect 301682 359360 301688 359372
rect 301280 359332 301688 359360
rect 301280 359320 301286 359332
rect 301682 359320 301688 359332
rect 301740 359360 301746 359372
rect 301792 359360 301820 359400
rect 306926 359388 306932 359400
rect 306984 359388 306990 359440
rect 307018 359388 307024 359440
rect 307076 359428 307082 359440
rect 312538 359428 312544 359440
rect 307076 359400 312544 359428
rect 307076 359388 307082 359400
rect 312538 359388 312544 359400
rect 312596 359388 312602 359440
rect 301740 359332 301820 359360
rect 301740 359320 301746 359332
rect 306926 359252 306932 359304
rect 306984 359292 306990 359304
rect 312262 359292 312268 359304
rect 306984 359264 312268 359292
rect 306984 359252 306990 359264
rect 312262 359252 312268 359264
rect 312320 359252 312326 359304
rect 273438 359184 273444 359236
rect 273496 359224 273502 359236
rect 278498 359224 278504 359236
rect 273496 359196 278504 359224
rect 273496 359184 273502 359196
rect 278498 359184 278504 359196
rect 278556 359184 278562 359236
rect 278590 359184 278596 359236
rect 278648 359224 278654 359236
rect 288802 359224 288808 359236
rect 278648 359196 288808 359224
rect 278648 359184 278654 359196
rect 288802 359184 288808 359196
rect 288860 359184 288866 359236
rect 292942 359184 292948 359236
rect 293000 359224 293006 359236
rect 294322 359224 294328 359236
rect 293000 359196 294328 359224
rect 293000 359184 293006 359196
rect 294322 359184 294328 359196
rect 294380 359224 294386 359236
rect 307018 359224 307024 359236
rect 294380 359196 307024 359224
rect 294380 359184 294386 359196
rect 307018 359184 307024 359196
rect 307076 359184 307082 359236
rect 307570 359184 307576 359236
rect 307628 359224 307634 359236
rect 312446 359224 312452 359236
rect 307628 359196 312452 359224
rect 307628 359184 307634 359196
rect 312446 359184 312452 359196
rect 312504 359184 312510 359236
rect 305270 358504 305276 358556
rect 305328 358544 305334 358556
rect 579246 358544 579252 358556
rect 305328 358516 579252 358544
rect 305328 358504 305334 358516
rect 579246 358504 579252 358516
rect 579304 358504 579310 358556
rect 267090 358436 267096 358488
rect 267148 358476 267154 358488
rect 294966 358476 294972 358488
rect 267148 358448 294972 358476
rect 267148 358436 267154 358448
rect 294966 358436 294972 358448
rect 295024 358436 295030 358488
rect 303246 358436 303252 358488
rect 303304 358476 303310 358488
rect 579338 358476 579344 358488
rect 303304 358448 579344 358476
rect 303304 358436 303310 358448
rect 579338 358436 579344 358448
rect 579396 358436 579402 358488
rect 3970 358368 3976 358420
rect 4028 358408 4034 358420
rect 274358 358408 274364 358420
rect 4028 358380 274364 358408
rect 4028 358368 4034 358380
rect 274358 358368 274364 358380
rect 274416 358368 274422 358420
rect 282638 358368 282644 358420
rect 282696 358408 282702 358420
rect 579614 358408 579620 358420
rect 282696 358380 579620 358408
rect 282696 358368 282702 358380
rect 579614 358368 579620 358380
rect 579672 358368 579678 358420
rect 299014 358300 299020 358352
rect 299072 358340 299078 358352
rect 300210 358340 300216 358352
rect 299072 358312 300216 358340
rect 299072 358300 299078 358312
rect 300210 358300 300216 358312
rect 300268 358300 300274 358352
rect 24946 357892 24952 357944
rect 25004 357932 25010 357944
rect 311342 357932 311348 357944
rect 25004 357904 311348 357932
rect 25004 357892 25010 357904
rect 311342 357892 311348 357904
rect 311400 357892 311406 357944
rect 271506 357824 271512 357876
rect 271564 357864 271570 357876
rect 296990 357864 296996 357876
rect 271564 357836 296996 357864
rect 271564 357824 271570 357836
rect 296990 357824 296996 357836
rect 297048 357824 297054 357876
rect 147122 357756 147128 357808
rect 147180 357796 147186 357808
rect 284662 357796 284668 357808
rect 147180 357768 284668 357796
rect 147180 357756 147186 357768
rect 284662 357756 284668 357768
rect 284720 357756 284726 357808
rect 290918 357756 290924 357808
rect 290976 357796 290982 357808
rect 317138 357796 317144 357808
rect 290976 357768 317144 357796
rect 290976 357756 290982 357768
rect 317138 357756 317144 357768
rect 317196 357756 317202 357808
rect 309318 357688 309324 357740
rect 309376 357728 309382 357740
rect 315666 357728 315672 357740
rect 309376 357700 315672 357728
rect 309376 357688 309382 357700
rect 315666 357688 315672 357700
rect 315724 357688 315730 357740
rect 273254 356260 273260 356312
rect 273312 356300 273318 356312
rect 275922 356300 275928 356312
rect 273312 356272 275928 356300
rect 273312 356260 273318 356272
rect 275922 356260 275928 356272
rect 275980 356260 275986 356312
rect 273530 354832 273536 354884
rect 273588 354872 273594 354884
rect 279694 354872 279700 354884
rect 273588 354844 279700 354872
rect 273588 354832 273594 354844
rect 279694 354832 279700 354844
rect 279752 354872 279758 354884
rect 280246 354872 280252 354884
rect 279752 354844 280252 354872
rect 279752 354832 279758 354844
rect 280246 354832 280252 354844
rect 280304 354832 280310 354884
rect 3878 354084 3884 354136
rect 3936 354124 3942 354136
rect 311526 354124 311532 354136
rect 3936 354096 311532 354124
rect 3936 354084 3942 354096
rect 311526 354084 311532 354096
rect 311584 354084 311590 354136
rect 270310 354016 270316 354068
rect 270368 354056 270374 354068
rect 579430 354056 579436 354068
rect 270368 354028 579436 354056
rect 270368 354016 270374 354028
rect 579430 354016 579436 354028
rect 579488 354016 579494 354068
rect 3786 353948 3792 354000
rect 3844 353988 3850 354000
rect 313550 353988 313556 354000
rect 3844 353960 313556 353988
rect 3844 353948 3850 353960
rect 313550 353948 313556 353960
rect 313608 353948 313614 354000
rect 269850 353200 269856 353252
rect 269908 353240 269914 353252
rect 270126 353240 270132 353252
rect 269908 353212 270132 353240
rect 269908 353200 269914 353212
rect 270126 353200 270132 353212
rect 270184 353200 270190 353252
rect 269666 350276 269672 350328
rect 269724 350316 269730 350328
rect 269850 350316 269856 350328
rect 269724 350288 269856 350316
rect 269724 350276 269730 350288
rect 269850 350276 269856 350288
rect 269908 350276 269914 350328
rect 269666 340076 269672 340128
rect 269724 340076 269730 340128
rect 269684 340048 269712 340076
rect 269942 340048 269948 340060
rect 269684 340020 269948 340048
rect 269942 340008 269948 340020
rect 270000 340008 270006 340060
rect 268562 339940 268568 339992
rect 268620 339980 268626 339992
rect 269666 339980 269672 339992
rect 268620 339952 269672 339980
rect 268620 339940 268626 339952
rect 269666 339940 269672 339952
rect 269724 339940 269730 339992
rect 314010 334092 314016 334144
rect 314068 334132 314074 334144
rect 579154 334132 579160 334144
rect 314068 334104 579160 334132
rect 314068 334092 314074 334104
rect 579154 334092 579160 334104
rect 579212 334092 579218 334144
rect 314010 333412 314016 333464
rect 314068 333452 314074 333464
rect 314286 333452 314292 333464
rect 314068 333424 314292 333452
rect 314068 333412 314074 333424
rect 314286 333412 314292 333424
rect 314344 333412 314350 333464
rect 268562 329740 268568 329792
rect 268620 329780 268626 329792
rect 269390 329780 269396 329792
rect 268620 329752 269396 329780
rect 268620 329740 268626 329752
rect 269390 329740 269396 329752
rect 269448 329740 269454 329792
rect 272150 316208 272156 316260
rect 272208 316248 272214 316260
rect 275278 316248 275284 316260
rect 272208 316220 275284 316248
rect 272208 316208 272214 316220
rect 275278 316208 275284 316220
rect 275336 316208 275342 316260
rect 310882 316208 310888 316260
rect 310940 316248 310946 316260
rect 312722 316248 312728 316260
rect 310940 316220 312728 316248
rect 310940 316208 310946 316220
rect 312722 316208 312728 316220
rect 312780 316208 312786 316260
rect 3602 313488 3608 313540
rect 3660 313528 3666 313540
rect 308582 313528 308588 313540
rect 3660 313500 308588 313528
rect 3660 313488 3666 313500
rect 308582 313488 308588 313500
rect 308640 313488 308646 313540
rect 3694 313420 3700 313472
rect 3752 313460 3758 313472
rect 285950 313460 285956 313472
rect 3752 313432 285956 313460
rect 3752 313420 3758 313432
rect 285950 313420 285956 313432
rect 286008 313420 286014 313472
rect 287974 313420 287980 313472
rect 288032 313460 288038 313472
rect 579522 313460 579528 313472
rect 288032 313432 579528 313460
rect 288032 313420 288038 313432
rect 579522 313420 579528 313432
rect 579580 313420 579586 313472
rect 272242 313352 272248 313404
rect 272300 313392 272306 313404
rect 283926 313392 283932 313404
rect 272300 313364 283932 313392
rect 272300 313352 272306 313364
rect 283926 313352 283932 313364
rect 283984 313352 283990 313404
rect 292206 313352 292212 313404
rect 292264 313392 292270 313404
rect 561490 313392 561496 313404
rect 292264 313364 561496 313392
rect 292264 313352 292270 313364
rect 561490 313352 561496 313364
rect 561548 313352 561554 313404
rect 24854 313284 24860 313336
rect 24912 313324 24918 313336
rect 273622 313324 273628 313336
rect 24912 313296 273628 313324
rect 24912 313284 24918 313296
rect 273622 313284 273628 313296
rect 273680 313284 273686 313336
rect 277670 313284 277676 313336
rect 277728 313324 277734 313336
rect 312814 313324 312820 313336
rect 277728 313296 312820 313324
rect 277728 313284 277734 313296
rect 312814 313284 312820 313296
rect 312872 313284 312878 313336
rect 271966 313216 271972 313268
rect 272024 313256 272030 313268
rect 281902 313256 281908 313268
rect 272024 313228 281908 313256
rect 272024 313216 272030 313228
rect 281902 313216 281908 313228
rect 281960 313216 281966 313268
rect 296254 313216 296260 313268
rect 296312 313256 296318 313268
rect 297266 313256 297272 313268
rect 296312 313228 297272 313256
rect 296312 313216 296318 313228
rect 297266 313216 297272 313228
rect 297324 313256 297330 313268
rect 313918 313256 313924 313268
rect 297324 313228 313924 313256
rect 297324 313216 297330 313228
rect 313918 313216 313924 313228
rect 313976 313216 313982 313268
rect 272058 313148 272064 313200
rect 272116 313188 272122 313200
rect 279694 313188 279700 313200
rect 272116 313160 279700 313188
rect 272116 313148 272122 313160
rect 279694 313148 279700 313160
rect 279752 313148 279758 313200
rect 298738 313148 298744 313200
rect 298796 313188 298802 313200
rect 313642 313188 313648 313200
rect 298796 313160 313648 313188
rect 298796 313148 298802 313160
rect 313642 313148 313648 313160
rect 313700 313148 313706 313200
rect 306558 313012 306564 313064
rect 306616 313052 306622 313064
rect 307570 313052 307576 313064
rect 306616 313024 307576 313052
rect 306616 313012 306622 313024
rect 307570 313012 307576 313024
rect 307628 313052 307634 313064
rect 313734 313052 313740 313064
rect 307628 313024 313740 313052
rect 307628 313012 307634 313024
rect 313734 313012 313740 313024
rect 313792 313012 313798 313064
rect 122098 312876 122104 312928
rect 122156 312916 122162 312928
rect 289998 312916 290004 312928
rect 122156 312888 290004 312916
rect 122156 312876 122162 312888
rect 289998 312876 290004 312888
rect 290056 312876 290062 312928
rect 98546 312808 98552 312860
rect 98604 312848 98610 312860
rect 300302 312848 300308 312860
rect 98604 312820 300308 312848
rect 98604 312808 98610 312820
rect 300302 312808 300308 312820
rect 300360 312808 300366 312860
rect 24854 312740 24860 312792
rect 24912 312780 24918 312792
rect 302510 312780 302516 312792
rect 24912 312752 302516 312780
rect 24912 312740 24918 312752
rect 302510 312740 302516 312752
rect 302568 312740 302574 312792
rect 270034 312128 270040 312180
rect 270092 312128 270098 312180
rect 270052 312044 270080 312128
rect 281166 312060 281172 312112
rect 281224 312100 281230 312112
rect 281902 312100 281908 312112
rect 281224 312072 281908 312100
rect 281224 312060 281230 312072
rect 281902 312060 281908 312072
rect 281960 312060 281966 312112
rect 282638 312060 282644 312112
rect 282696 312100 282702 312112
rect 283926 312100 283932 312112
rect 282696 312072 283932 312100
rect 282696 312060 282702 312072
rect 283926 312060 283932 312072
rect 283984 312060 283990 312112
rect 270034 311992 270040 312044
rect 270092 311992 270098 312044
rect 303890 311992 303896 312044
rect 303948 312032 303954 312044
rect 304534 312032 304540 312044
rect 303948 312004 304540 312032
rect 303948 311992 303954 312004
rect 304534 311992 304540 312004
rect 304592 312032 304598 312044
rect 312630 312032 312636 312044
rect 304592 312004 312636 312032
rect 304592 311992 304598 312004
rect 312630 311992 312636 312004
rect 312688 311992 312694 312044
rect 270034 309068 270040 309120
rect 270092 309108 270098 309120
rect 270310 309108 270316 309120
rect 270092 309080 270316 309108
rect 270092 309068 270098 309080
rect 270310 309068 270316 309080
rect 270368 309068 270374 309120
rect 269850 291456 269856 291508
rect 269908 291456 269914 291508
rect 269868 291360 269896 291456
rect 269942 291360 269948 291372
rect 269868 291332 269948 291360
rect 269942 291320 269948 291332
rect 270000 291320 270006 291372
rect 97994 276700 98000 276752
rect 98052 276740 98058 276752
rect 98546 276740 98552 276752
rect 98052 276712 98552 276740
rect 98052 276700 98058 276712
rect 98546 276700 98552 276712
rect 98604 276700 98610 276752
rect 146202 276700 146208 276752
rect 146260 276740 146266 276752
rect 147122 276740 147128 276752
rect 146260 276712 147128 276740
rect 146260 276700 146266 276712
rect 147122 276700 147128 276712
rect 147180 276700 147186 276752
rect 170122 276632 170128 276684
rect 170180 276672 170186 276684
rect 175182 276672 175188 276684
rect 170180 276644 175188 276672
rect 170180 276632 170186 276644
rect 175182 276632 175188 276644
rect 175240 276632 175246 276684
rect 195790 276672 195796 276684
rect 190564 276644 195796 276672
rect 185394 276564 185400 276616
rect 185452 276604 185458 276616
rect 188338 276604 188344 276616
rect 185452 276576 188344 276604
rect 185452 276564 185458 276576
rect 188338 276564 188344 276576
rect 188396 276564 188402 276616
rect 188430 276564 188436 276616
rect 188488 276604 188494 276616
rect 190564 276604 190592 276644
rect 195790 276632 195796 276644
rect 195848 276632 195854 276684
rect 216398 276672 216404 276684
rect 211172 276644 216404 276672
rect 188488 276576 190592 276604
rect 188488 276564 188494 276576
rect 206002 276564 206008 276616
rect 206060 276604 206066 276616
rect 208946 276604 208952 276616
rect 206060 276576 208952 276604
rect 206060 276564 206066 276576
rect 208946 276564 208952 276576
rect 209004 276564 209010 276616
rect 209038 276564 209044 276616
rect 209096 276604 209102 276616
rect 211172 276604 211200 276644
rect 216398 276632 216404 276644
rect 216456 276632 216462 276684
rect 237006 276672 237012 276684
rect 231780 276644 237012 276672
rect 209096 276576 211200 276604
rect 209096 276564 209102 276576
rect 226610 276564 226616 276616
rect 226668 276604 226674 276616
rect 229554 276604 229560 276616
rect 226668 276576 229560 276604
rect 226668 276564 226674 276576
rect 229554 276564 229560 276576
rect 229612 276564 229618 276616
rect 229646 276564 229652 276616
rect 229704 276604 229710 276616
rect 231780 276604 231808 276644
rect 237006 276632 237012 276644
rect 237064 276632 237070 276684
rect 257614 276632 257620 276684
rect 257672 276672 257678 276684
rect 267826 276672 267832 276684
rect 257672 276644 267832 276672
rect 257672 276632 257678 276644
rect 267826 276632 267832 276644
rect 267884 276632 267890 276684
rect 229704 276576 231808 276604
rect 229704 276564 229710 276576
rect 240042 276564 240048 276616
rect 240100 276604 240106 276616
rect 250254 276604 250260 276616
rect 240100 276576 250260 276604
rect 240100 276564 240106 276576
rect 250254 276564 250260 276576
rect 250312 276564 250318 276616
rect 285582 276564 285588 276616
rect 285640 276604 285646 276616
rect 295794 276604 295800 276616
rect 285640 276576 295800 276604
rect 285640 276564 285646 276576
rect 295794 276564 295800 276576
rect 295852 276564 295858 276616
rect 307018 276564 307024 276616
rect 307076 276604 307082 276616
rect 307570 276604 307576 276616
rect 307076 276576 307576 276604
rect 307076 276564 307082 276576
rect 307570 276564 307576 276576
rect 307628 276604 307634 276616
rect 341794 276604 341800 276616
rect 307628 276576 341800 276604
rect 307628 276564 307634 276576
rect 341794 276564 341800 276576
rect 341852 276564 341858 276616
rect 242434 276496 242440 276548
rect 242492 276536 242498 276548
rect 312078 276536 312084 276548
rect 242492 276508 312084 276536
rect 242492 276496 242498 276508
rect 312078 276496 312084 276508
rect 312136 276536 312142 276548
rect 312538 276536 312544 276548
rect 312136 276508 312544 276536
rect 312136 276496 312142 276508
rect 312538 276496 312544 276508
rect 312596 276496 312602 276548
rect 326890 276496 326896 276548
rect 326948 276536 326954 276548
rect 337010 276536 337016 276548
rect 326948 276508 337016 276536
rect 326948 276496 326954 276508
rect 337010 276496 337016 276508
rect 337068 276496 337074 276548
rect 347498 276496 347504 276548
rect 347556 276536 347562 276548
rect 357618 276536 357624 276548
rect 347556 276508 357624 276536
rect 347556 276496 347562 276508
rect 357618 276496 357624 276508
rect 357676 276496 357682 276548
rect 365714 276536 365720 276548
rect 359200 276508 365720 276536
rect 257614 276428 257620 276480
rect 257672 276428 257678 276480
rect 267826 276428 267832 276480
rect 267884 276468 267890 276480
rect 267884 276440 270908 276468
rect 267884 276428 267890 276440
rect 250254 276360 250260 276412
rect 250312 276400 250318 276412
rect 257632 276400 257660 276428
rect 250312 276372 257660 276400
rect 270880 276400 270908 276440
rect 282638 276428 282644 276480
rect 282696 276468 282702 276480
rect 359200 276468 359228 276508
rect 365714 276496 365720 276508
rect 365772 276496 365778 276548
rect 403986 276496 403992 276548
rect 404044 276536 404050 276548
rect 419442 276536 419448 276548
rect 404044 276508 419448 276536
rect 404044 276496 404050 276508
rect 419442 276496 419448 276508
rect 419500 276496 419506 276548
rect 443086 276536 443092 276548
rect 437860 276508 443092 276536
rect 282696 276440 359228 276468
rect 282696 276428 282702 276440
rect 362770 276428 362776 276480
rect 362828 276468 362834 276480
rect 378226 276468 378232 276480
rect 362828 276440 378232 276468
rect 362828 276428 362834 276440
rect 378226 276428 378232 276440
rect 378284 276428 378290 276480
rect 383378 276428 383384 276480
rect 383436 276468 383442 276480
rect 398834 276468 398840 276480
rect 383436 276440 398840 276468
rect 383436 276428 383442 276440
rect 398834 276428 398840 276440
rect 398892 276428 398898 276480
rect 429838 276428 429844 276480
rect 429896 276468 429902 276480
rect 435634 276468 435640 276480
rect 429896 276440 435640 276468
rect 429896 276428 429902 276440
rect 435634 276428 435640 276440
rect 435692 276428 435698 276480
rect 435726 276428 435732 276480
rect 435784 276468 435790 276480
rect 437860 276468 437888 276508
rect 443086 276496 443092 276508
rect 443144 276496 443150 276548
rect 435784 276440 437888 276468
rect 435784 276428 435790 276440
rect 453298 276428 453304 276480
rect 453356 276468 453362 276480
rect 454218 276468 454224 276480
rect 453356 276440 454224 276468
rect 453356 276428 453362 276440
rect 454218 276428 454224 276440
rect 454276 276428 454282 276480
rect 270880 276372 281120 276400
rect 250312 276360 250318 276372
rect 281092 276332 281120 276372
rect 294322 276360 294328 276412
rect 294380 276400 294386 276412
rect 413922 276400 413928 276412
rect 294380 276372 413928 276400
rect 294380 276360 294386 276372
rect 413922 276360 413928 276372
rect 413980 276360 413986 276412
rect 285582 276332 285588 276344
rect 281092 276304 285588 276332
rect 285582 276292 285588 276304
rect 285640 276292 285646 276344
rect 317138 276292 317144 276344
rect 317196 276332 317202 276344
rect 438026 276332 438032 276344
rect 317196 276304 438032 276332
rect 317196 276292 317202 276304
rect 438026 276292 438032 276304
rect 438084 276292 438090 276344
rect 73522 276224 73528 276276
rect 73580 276264 73586 276276
rect 282638 276264 282644 276276
rect 73580 276236 282644 276264
rect 73580 276224 73586 276236
rect 282638 276224 282644 276236
rect 282696 276224 282702 276276
rect 295794 276224 295800 276276
rect 295852 276264 295858 276276
rect 298738 276264 298744 276276
rect 295852 276236 298744 276264
rect 295852 276224 295858 276236
rect 298738 276224 298744 276236
rect 298796 276264 298802 276276
rect 306190 276264 306196 276276
rect 298796 276236 306196 276264
rect 298796 276224 298802 276236
rect 306190 276224 306196 276236
rect 306248 276224 306254 276276
rect 316402 276224 316408 276276
rect 316460 276264 316466 276276
rect 326890 276264 326896 276276
rect 316460 276236 326896 276264
rect 316460 276224 316466 276236
rect 326890 276224 326896 276236
rect 326948 276224 326954 276276
rect 337010 276224 337016 276276
rect 337068 276264 337074 276276
rect 347498 276264 347504 276276
rect 337068 276236 347504 276264
rect 337068 276224 337074 276236
rect 347498 276224 347504 276236
rect 347556 276224 347562 276276
rect 357618 276224 357624 276276
rect 357676 276264 357682 276276
rect 362770 276264 362776 276276
rect 357676 276236 362776 276264
rect 357676 276224 357682 276236
rect 362770 276224 362776 276236
rect 362828 276224 362834 276276
rect 378226 276224 378232 276276
rect 378284 276264 378290 276276
rect 383378 276264 383384 276276
rect 378284 276236 383384 276264
rect 378284 276224 378290 276236
rect 383378 276224 383384 276236
rect 383436 276224 383442 276276
rect 398834 276224 398840 276276
rect 398892 276264 398898 276276
rect 403986 276264 403992 276276
rect 398892 276236 403992 276264
rect 398892 276224 398898 276236
rect 403986 276224 403992 276236
rect 404044 276224 404050 276276
rect 419442 276224 419448 276276
rect 419500 276264 419506 276276
rect 429838 276264 429844 276276
rect 419500 276236 429844 276264
rect 419500 276224 419506 276236
rect 429838 276224 429844 276236
rect 429896 276224 429902 276276
rect 454218 276224 454224 276276
rect 454276 276264 454282 276276
rect 461946 276264 461952 276276
rect 454276 276236 461952 276264
rect 454276 276224 454282 276236
rect 461946 276224 461952 276236
rect 462004 276224 462010 276276
rect 194226 276156 194232 276208
rect 194284 276196 194290 276208
rect 270402 276196 270408 276208
rect 194284 276168 270408 276196
rect 194284 276156 194290 276168
rect 270402 276156 270408 276168
rect 270460 276196 270466 276208
rect 486050 276196 486056 276208
rect 270460 276168 486056 276196
rect 270460 276156 270466 276168
rect 486050 276156 486056 276168
rect 486108 276156 486114 276208
rect 218330 276088 218336 276140
rect 218388 276128 218394 276140
rect 270218 276128 270224 276140
rect 218388 276100 270224 276128
rect 218388 276088 218394 276100
rect 270218 276088 270224 276100
rect 270276 276128 270282 276140
rect 510154 276128 510160 276140
rect 270276 276100 510160 276128
rect 270276 276088 270282 276100
rect 510154 276088 510160 276100
rect 510212 276088 510218 276140
rect 49970 276020 49976 276072
rect 50028 276060 50034 276072
rect 307018 276060 307024 276072
rect 50028 276032 307024 276060
rect 50028 276020 50034 276032
rect 307018 276020 307024 276032
rect 307076 276020 307082 276072
rect 312078 276020 312084 276072
rect 312136 276060 312142 276072
rect 534258 276060 534264 276072
rect 312136 276032 534264 276060
rect 312136 276020 312142 276032
rect 534258 276020 534264 276032
rect 534316 276020 534322 276072
rect 266354 275952 266360 276004
rect 266412 275992 266418 276004
rect 273162 275992 273168 276004
rect 266412 275964 273168 275992
rect 266412 275952 266418 275964
rect 273162 275952 273168 275964
rect 273220 275992 273226 276004
rect 558178 275992 558184 276004
rect 273220 275964 558184 275992
rect 273220 275952 273226 275964
rect 558178 275952 558184 275964
rect 558236 275952 558242 276004
rect 306190 275884 306196 275936
rect 306248 275924 306254 275936
rect 316402 275924 316408 275936
rect 306248 275896 316408 275924
rect 306248 275884 306254 275896
rect 316402 275884 316408 275896
rect 316460 275884 316466 275936
rect 314378 272348 314384 272400
rect 314436 272388 314442 272400
rect 560846 272388 560852 272400
rect 314436 272360 560852 272388
rect 314436 272348 314442 272360
rect 560846 272348 560852 272360
rect 560904 272348 560910 272400
rect 275922 272212 275928 272264
rect 275980 272252 275986 272264
rect 275980 272224 285536 272252
rect 275980 272212 275986 272224
rect 26418 272076 26424 272128
rect 26476 272116 26482 272128
rect 273254 272116 273260 272128
rect 26476 272088 273260 272116
rect 26476 272076 26482 272088
rect 273254 272076 273260 272088
rect 273312 272116 273318 272128
rect 276658 272116 276664 272128
rect 273312 272088 276664 272116
rect 273312 272076 273318 272088
rect 276658 272076 276664 272088
rect 276716 272076 276722 272128
rect 285508 272116 285536 272224
rect 558638 272116 558644 272128
rect 285508 272088 558644 272116
rect 558638 272076 558644 272088
rect 558696 272076 558702 272128
rect 27154 272008 27160 272060
rect 27212 272048 27218 272060
rect 312538 272048 312544 272060
rect 27212 272020 312544 272048
rect 27212 272008 27218 272020
rect 312538 272008 312544 272020
rect 312596 272008 312602 272060
rect 27614 271940 27620 271992
rect 27672 271980 27678 271992
rect 314010 271980 314016 271992
rect 27672 271952 314016 271980
rect 27672 271940 27678 271952
rect 314010 271940 314016 271952
rect 314068 271940 314074 271992
rect 314010 270852 314016 270904
rect 314068 270892 314074 270904
rect 314286 270892 314292 270904
rect 314068 270864 314292 270892
rect 314068 270852 314074 270864
rect 314286 270852 314292 270864
rect 314344 270852 314350 270904
rect 276658 270784 276664 270836
rect 276716 270824 276722 270836
rect 315022 270824 315028 270836
rect 276716 270796 315028 270824
rect 276716 270784 276722 270796
rect 315022 270784 315028 270796
rect 315080 270784 315086 270836
rect 26142 267928 26148 267980
rect 26200 267968 26206 267980
rect 27614 267968 27620 267980
rect 26200 267940 27620 267968
rect 26200 267928 26206 267940
rect 27614 267928 27620 267940
rect 27672 267928 27678 267980
rect 558454 267928 558460 267980
rect 558512 267968 558518 267980
rect 558638 267968 558644 267980
rect 558512 267940 558644 267968
rect 558512 267928 558518 267940
rect 558638 267928 558644 267940
rect 558696 267928 558702 267980
rect 558546 257524 558552 257576
rect 558604 257564 558610 257576
rect 558638 257564 558644 257576
rect 558604 257536 558644 257564
rect 558604 257524 558610 257536
rect 558638 257524 558644 257536
rect 558696 257524 558702 257576
rect 24762 256164 24768 256216
rect 24820 256204 24826 256216
rect 27154 256204 27160 256216
rect 24820 256176 27160 256204
rect 24820 256164 24826 256176
rect 27154 256164 27160 256176
rect 27212 256164 27218 256216
rect 558546 247256 558552 247308
rect 558604 247296 558610 247308
rect 558730 247296 558736 247308
rect 558604 247268 558736 247296
rect 558604 247256 558610 247268
rect 558730 247256 558736 247268
rect 558788 247256 558794 247308
rect 268378 238416 268384 238468
rect 268436 238456 268442 238468
rect 314378 238456 314384 238468
rect 268436 238428 314384 238456
rect 268436 238416 268442 238428
rect 314378 238416 314384 238428
rect 314436 238416 314442 238468
rect 270126 236988 270132 237040
rect 270184 237028 270190 237040
rect 270218 237028 270224 237040
rect 270184 237000 270224 237028
rect 270184 236988 270190 237000
rect 270218 236988 270224 237000
rect 270276 236988 270282 237040
rect 558546 236988 558552 237040
rect 558604 237028 558610 237040
rect 558822 237028 558828 237040
rect 558604 237000 558828 237028
rect 558604 236988 558610 237000
rect 558822 236988 558828 237000
rect 558880 236988 558886 237040
rect 558822 229752 558828 229764
rect 558748 229724 558828 229752
rect 558748 229628 558776 229724
rect 558822 229712 558828 229724
rect 558880 229712 558886 229764
rect 558730 229576 558736 229628
rect 558788 229576 558794 229628
rect 269850 226720 269856 226772
rect 269908 226760 269914 226772
rect 270218 226760 270224 226772
rect 269908 226732 270224 226760
rect 269908 226720 269914 226732
rect 270218 226720 270224 226732
rect 270276 226720 270282 226772
rect 270126 216384 270132 216436
rect 270184 216424 270190 216436
rect 270218 216424 270224 216436
rect 270184 216396 270224 216424
rect 270184 216384 270190 216396
rect 270218 216384 270224 216396
rect 270276 216384 270282 216436
rect 270218 206048 270224 206100
rect 270276 206088 270282 206100
rect 270402 206088 270408 206100
rect 270276 206060 270408 206088
rect 270276 206048 270282 206060
rect 270402 206048 270408 206060
rect 270460 206048 270466 206100
rect 558454 203124 558460 203176
rect 558512 203164 558518 203176
rect 558822 203164 558828 203176
rect 558512 203136 558828 203164
rect 558512 203124 558518 203136
rect 558822 203124 558828 203136
rect 558880 203124 558886 203176
rect 268378 202784 268384 202836
rect 268436 202824 268442 202836
rect 275922 202824 275928 202836
rect 268436 202796 275928 202824
rect 268436 202784 268442 202796
rect 275922 202784 275928 202796
rect 275980 202784 275986 202836
rect 312722 200132 312728 200184
rect 312780 200172 312786 200184
rect 315022 200172 315028 200184
rect 312780 200144 315028 200172
rect 312780 200132 312786 200144
rect 315022 200132 315028 200144
rect 315080 200132 315086 200184
rect 270126 195780 270132 195832
rect 270184 195820 270190 195832
rect 270402 195820 270408 195832
rect 270184 195792 270408 195820
rect 270184 195780 270190 195792
rect 270402 195780 270408 195792
rect 270460 195780 270466 195832
rect 270218 185444 270224 185496
rect 270276 185484 270282 185496
rect 270402 185484 270408 185496
rect 270276 185456 270408 185484
rect 270276 185444 270282 185456
rect 270402 185444 270408 185456
rect 270460 185444 270466 185496
rect 270126 175176 270132 175228
rect 270184 175216 270190 175228
rect 270402 175216 270408 175228
rect 270184 175188 270408 175216
rect 270184 175176 270190 175188
rect 270402 175176 270408 175188
rect 270460 175176 270466 175228
rect 270218 164772 270224 164824
rect 270276 164812 270282 164824
rect 270402 164812 270408 164824
rect 270276 164784 270408 164812
rect 270276 164772 270282 164784
rect 270402 164772 270408 164784
rect 270460 164772 270466 164824
rect 270126 147296 270132 147348
rect 270184 147296 270190 147348
rect 270144 147212 270172 147296
rect 270126 147160 270132 147212
rect 270184 147160 270190 147212
rect 270126 144236 270132 144288
rect 270184 144276 270190 144288
rect 270218 144276 270224 144288
rect 270184 144248 270224 144276
rect 270184 144236 270190 144248
rect 270218 144236 270224 144248
rect 270276 144236 270282 144288
rect 270126 142740 270132 142792
rect 270184 142780 270190 142792
rect 270402 142780 270408 142792
rect 270184 142752 270408 142780
rect 270184 142740 270190 142752
rect 270402 142740 270408 142752
rect 270460 142740 270466 142792
rect 270126 132472 270132 132524
rect 270184 132472 270190 132524
rect 270144 132444 270172 132472
rect 270218 132444 270224 132456
rect 270144 132416 270224 132444
rect 270218 132404 270224 132416
rect 270276 132404 270282 132456
rect 268286 130568 268292 130620
rect 268344 130608 268350 130620
rect 273346 130608 273352 130620
rect 268344 130580 273352 130608
rect 268344 130568 268350 130580
rect 273346 130568 273352 130580
rect 273404 130568 273410 130620
rect 273346 130228 273352 130280
rect 273404 130268 273410 130280
rect 291470 130268 291476 130280
rect 273404 130240 291476 130268
rect 273404 130228 273410 130240
rect 291470 130228 291476 130240
rect 291528 130228 291534 130280
rect 270126 126624 270132 126676
rect 270184 126624 270190 126676
rect 270144 126528 270172 126624
rect 270218 126528 270224 126540
rect 270144 126500 270224 126528
rect 270218 126488 270224 126500
rect 270276 126488 270282 126540
rect 558546 125604 558552 125656
rect 558604 125644 558610 125656
rect 559374 125644 559380 125656
rect 558604 125616 559380 125644
rect 558604 125604 558610 125616
rect 559374 125604 559380 125616
rect 559432 125604 559438 125656
rect 291470 125536 291476 125588
rect 291528 125576 291534 125588
rect 293586 125576 293592 125588
rect 291528 125548 293592 125576
rect 291528 125536 291534 125548
rect 293586 125536 293592 125548
rect 293644 125536 293650 125588
rect 270218 116288 270224 116340
rect 270276 116288 270282 116340
rect 270236 116192 270264 116288
rect 293586 116220 293592 116272
rect 293644 116260 293650 116272
rect 294690 116260 294696 116272
rect 293644 116232 294696 116260
rect 293644 116220 293650 116232
rect 294690 116220 294696 116232
rect 294748 116220 294754 116272
rect 270310 116192 270316 116204
rect 270236 116164 270316 116192
rect 270310 116152 270316 116164
rect 270368 116152 270374 116204
rect 294690 114724 294696 114776
rect 294748 114764 294754 114776
rect 296438 114764 296444 114776
rect 294748 114736 296444 114764
rect 294748 114724 294754 114736
rect 296438 114724 296444 114736
rect 296496 114724 296502 114776
rect 296438 111800 296444 111852
rect 296496 111840 296502 111852
rect 297358 111840 297364 111852
rect 296496 111812 297364 111840
rect 296496 111800 296502 111812
rect 297358 111800 297364 111812
rect 297416 111800 297422 111852
rect 297358 109284 297364 109336
rect 297416 109324 297422 109336
rect 300210 109324 300216 109336
rect 297416 109296 300216 109324
rect 297416 109284 297422 109296
rect 300210 109284 300216 109296
rect 300268 109284 300274 109336
rect 270218 101600 270224 101652
rect 270276 101640 270282 101652
rect 270310 101640 270316 101652
rect 270276 101612 270316 101640
rect 270276 101600 270282 101612
rect 270310 101600 270316 101612
rect 270368 101600 270374 101652
rect 300302 101532 300308 101584
rect 300360 101572 300366 101584
rect 301774 101572 301780 101584
rect 300360 101544 301780 101572
rect 300360 101532 300366 101544
rect 301774 101532 301780 101544
rect 301832 101532 301838 101584
rect 267918 94868 267924 94920
rect 267976 94908 267982 94920
rect 303890 94908 303896 94920
rect 267976 94880 303896 94908
rect 267976 94868 267982 94880
rect 303890 94868 303896 94880
rect 303948 94868 303954 94920
rect 301774 94188 301780 94240
rect 301832 94228 301838 94240
rect 301832 94200 303292 94228
rect 301832 94188 301838 94200
rect 303264 94160 303292 94200
rect 304718 94160 304724 94172
rect 303264 94132 304724 94160
rect 304718 94120 304724 94132
rect 304776 94120 304782 94172
rect 314194 92352 314200 92404
rect 314252 92392 314258 92404
rect 315022 92392 315028 92404
rect 314252 92364 315028 92392
rect 314252 92352 314258 92364
rect 315022 92352 315028 92364
rect 315080 92352 315086 92404
rect 269942 91264 269948 91316
rect 270000 91304 270006 91316
rect 270126 91304 270132 91316
rect 270000 91276 270132 91304
rect 270000 91264 270006 91276
rect 270126 91264 270132 91276
rect 270184 91264 270190 91316
rect 304718 90380 304724 90432
rect 304776 90420 304782 90432
rect 307662 90420 307668 90432
rect 304776 90392 307668 90420
rect 304776 90380 304782 90392
rect 307662 90380 307668 90392
rect 307720 90380 307726 90432
rect 307662 86844 307668 86896
rect 307720 86884 307726 86896
rect 307720 86856 309180 86884
rect 307720 86844 307726 86856
rect 309152 86816 309180 86856
rect 312078 86816 312084 86828
rect 309152 86788 312084 86816
rect 312078 86776 312084 86788
rect 312136 86776 312142 86828
rect 269942 82424 269948 82476
rect 270000 82464 270006 82476
rect 270310 82464 270316 82476
rect 270000 82436 270316 82464
rect 270000 82424 270006 82436
rect 270310 82424 270316 82436
rect 270368 82424 270374 82476
rect 312078 81132 312084 81184
rect 312136 81172 312142 81184
rect 316494 81172 316500 81184
rect 312136 81144 316500 81172
rect 312136 81132 312142 81144
rect 316494 81132 316500 81144
rect 316552 81132 316558 81184
rect 24946 75964 24952 76016
rect 25004 76004 25010 76016
rect 314194 76004 314200 76016
rect 25004 75976 314200 76004
rect 25004 75964 25010 75976
rect 314194 75964 314200 75976
rect 314252 75964 314258 76016
rect 316494 75964 316500 76016
rect 316552 76004 316558 76016
rect 558546 76004 558552 76016
rect 316552 75976 558552 76004
rect 316552 75964 316558 75976
rect 558546 75964 558552 75976
rect 558604 75964 558610 76016
rect 303890 75896 303896 75948
rect 303948 75936 303954 75948
rect 560846 75936 560852 75948
rect 303948 75908 560852 75936
rect 303948 75896 303954 75908
rect 560846 75896 560852 75908
rect 560904 75896 560910 75948
rect 39666 72088 39672 72140
rect 39724 72128 39730 72140
rect 312354 72128 312360 72140
rect 39724 72100 312360 72128
rect 39724 72088 39730 72100
rect 312354 72088 312360 72100
rect 312412 72088 312418 72140
rect 313550 72088 313556 72140
rect 313608 72128 313614 72140
rect 475930 72128 475936 72140
rect 313608 72100 475936 72128
rect 313608 72088 313614 72100
rect 475930 72088 475936 72100
rect 475988 72088 475994 72140
rect 63770 72020 63776 72072
rect 63828 72060 63834 72072
rect 269390 72060 269396 72072
rect 63828 72032 269396 72060
rect 63828 72020 63834 72032
rect 269390 72020 269396 72032
rect 269448 72020 269454 72072
rect 279694 72020 279700 72072
rect 279752 72060 279758 72072
rect 280154 72060 280160 72072
rect 279752 72032 280160 72060
rect 279752 72020 279758 72032
rect 280154 72020 280160 72032
rect 280212 72060 280218 72072
rect 548058 72060 548064 72072
rect 280212 72032 548064 72060
rect 280212 72020 280218 72032
rect 548058 72020 548064 72032
rect 548116 72020 548122 72072
rect 272334 71952 272340 72004
rect 272392 71992 272398 72004
rect 273438 71992 273444 72004
rect 272392 71964 273444 71992
rect 272392 71952 272398 71964
rect 273438 71952 273444 71964
rect 273496 71992 273502 72004
rect 499850 71992 499856 72004
rect 273496 71964 499856 71992
rect 273496 71952 273502 71964
rect 499850 71952 499856 71964
rect 499908 71952 499914 72004
rect 87690 71884 87696 71936
rect 87748 71924 87754 71936
rect 281166 71924 281172 71936
rect 87748 71896 281172 71924
rect 87748 71884 87754 71896
rect 281166 71884 281172 71896
rect 281224 71884 281230 71936
rect 297266 71884 297272 71936
rect 297324 71924 297330 71936
rect 523954 71924 523960 71936
rect 297324 71896 523960 71924
rect 297324 71884 297330 71896
rect 523954 71884 523960 71896
rect 524012 71884 524018 71936
rect 135898 71816 135904 71868
rect 135956 71856 135962 71868
rect 314102 71856 314108 71868
rect 135956 71828 314108 71856
rect 135956 71816 135962 71828
rect 314102 71816 314108 71828
rect 314160 71856 314166 71868
rect 427722 71856 427728 71868
rect 314160 71828 427728 71856
rect 314160 71816 314166 71828
rect 427722 71816 427728 71828
rect 427780 71816 427786 71868
rect 183922 71748 183928 71800
rect 183980 71788 183986 71800
rect 313550 71788 313556 71800
rect 183980 71760 313556 71788
rect 183980 71748 183986 71760
rect 313550 71748 313556 71760
rect 313608 71748 313614 71800
rect 160002 71680 160008 71732
rect 160060 71720 160066 71732
rect 271506 71720 271512 71732
rect 160060 71692 271512 71720
rect 160060 71680 160066 71692
rect 271506 71680 271512 71692
rect 271564 71680 271570 71732
rect 272426 71680 272432 71732
rect 272484 71720 272490 71732
rect 273530 71720 273536 71732
rect 272484 71692 273536 71720
rect 272484 71680 272490 71692
rect 273530 71680 273536 71692
rect 273588 71720 273594 71732
rect 403618 71720 403624 71732
rect 273588 71692 403624 71720
rect 273588 71680 273594 71692
rect 403618 71680 403624 71692
rect 403676 71680 403682 71732
rect 208026 71612 208032 71664
rect 208084 71652 208090 71664
rect 272334 71652 272340 71664
rect 208084 71624 272340 71652
rect 208084 71612 208090 71624
rect 272334 71612 272340 71624
rect 272392 71612 272398 71664
rect 281166 71612 281172 71664
rect 281224 71652 281230 71664
rect 379514 71652 379520 71664
rect 281224 71624 379520 71652
rect 281224 71612 281230 71624
rect 379514 71612 379520 71624
rect 379572 71612 379578 71664
rect 269390 71544 269396 71596
rect 269448 71584 269454 71596
rect 270310 71584 270316 71596
rect 269448 71556 270316 71584
rect 269448 71544 269454 71556
rect 270310 71544 270316 71556
rect 270368 71584 270374 71596
rect 355594 71584 355600 71596
rect 270368 71556 355600 71584
rect 270368 71544 270374 71556
rect 355594 71544 355600 71556
rect 355652 71544 355658 71596
rect 232130 71476 232136 71528
rect 232188 71516 232194 71528
rect 297266 71516 297272 71528
rect 232188 71488 297272 71516
rect 232188 71476 232194 71488
rect 297266 71476 297272 71488
rect 297324 71476 297330 71528
rect 312354 71476 312360 71528
rect 312412 71516 312418 71528
rect 331490 71516 331496 71528
rect 312412 71488 331496 71516
rect 312412 71476 312418 71488
rect 331490 71476 331496 71488
rect 331548 71476 331554 71528
rect 256050 71408 256056 71460
rect 256108 71448 256114 71460
rect 280154 71448 280160 71460
rect 256108 71420 280160 71448
rect 256108 71408 256114 71420
rect 280154 71408 280160 71420
rect 280212 71408 280218 71460
rect 111794 71340 111800 71392
rect 111852 71380 111858 71392
rect 272426 71380 272432 71392
rect 111852 71352 272432 71380
rect 111852 71340 111858 71352
rect 272426 71340 272432 71352
rect 272484 71340 272490 71392
rect 270586 3612 270592 3664
rect 270644 3652 270650 3664
rect 583386 3652 583392 3664
rect 270644 3624 583392 3652
rect 270644 3612 270650 3624
rect 583386 3612 583392 3624
rect 583444 3612 583450 3664
<< via1 >>
rect 8024 700612 8076 700664
rect 8208 700612 8260 700664
rect 72976 700612 73028 700664
rect 137836 700612 137888 700664
rect 202788 700612 202840 700664
rect 267648 700612 267700 700664
rect 332508 700612 332560 700664
rect 397460 700612 397512 700664
rect 462320 700612 462372 700664
rect 527180 700612 527232 700664
rect 272984 700272 273036 700324
rect 283840 700272 283892 700324
rect 270868 700204 270920 700256
rect 364984 700204 365036 700256
rect 218980 700136 219032 700188
rect 312084 700136 312136 700188
rect 270684 700068 270736 700120
rect 429844 700068 429896 700120
rect 89168 700000 89220 700052
rect 312176 700000 312228 700052
rect 312728 700000 312780 700052
rect 494796 700000 494848 700052
rect 154120 699932 154172 699984
rect 268568 699932 268620 699984
rect 270776 699932 270828 699984
rect 559656 699932 559708 699984
rect 24308 699864 24360 699916
rect 314476 699864 314528 699916
rect 527180 699864 527232 699916
rect 579896 699864 579948 699916
rect 561496 674160 561548 674212
rect 578516 674160 578568 674212
rect 2964 653488 3016 653540
rect 8024 653488 8076 653540
rect 270500 627104 270552 627156
rect 578792 627104 578844 627156
rect 49608 586576 49660 586628
rect 313740 586576 313792 586628
rect 217968 586508 218020 586560
rect 270592 586508 270644 586560
rect 271144 586508 271196 586560
rect 306196 586508 306248 586560
rect 316408 586508 316460 586560
rect 326896 586508 326948 586560
rect 337016 586508 337068 586560
rect 347412 586508 347464 586560
rect 357624 586508 357676 586560
rect 73528 586440 73580 586492
rect 272248 586440 272300 586492
rect 365444 586440 365496 586492
rect 368020 586440 368072 586492
rect 378232 586440 378284 586492
rect 388628 586440 388680 586492
rect 398840 586440 398892 586492
rect 409236 586440 409288 586492
rect 415124 586440 415176 586492
rect 242072 586372 242124 586424
rect 292948 586372 293000 586424
rect 300216 586372 300268 586424
rect 437756 586372 437808 586424
rect 169760 586304 169812 586356
rect 313648 586304 313700 586356
rect 313740 586304 313792 586356
rect 341524 586304 341576 586356
rect 121736 586236 121788 586288
rect 312360 586236 312412 586288
rect 312820 586236 312872 586288
rect 413652 586236 413704 586288
rect 415124 586236 415176 586288
rect 198740 586168 198792 586220
rect 209044 586168 209096 586220
rect 216496 586168 216548 586220
rect 229652 586168 229704 586220
rect 239956 586100 240008 586152
rect 250260 586100 250312 586152
rect 145840 586032 145892 586084
rect 267096 586032 267148 586084
rect 193864 585964 193916 586016
rect 198740 585964 198792 586016
rect 229652 585964 229704 586016
rect 209044 585896 209096 585948
rect 216404 585896 216456 585948
rect 257620 585964 257672 586016
rect 267740 585964 267792 586016
rect 270408 586100 270460 586152
rect 306196 586168 306248 586220
rect 316408 586168 316460 586220
rect 326896 586168 326948 586220
rect 337016 586168 337068 586220
rect 347412 586168 347464 586220
rect 357624 586168 357676 586220
rect 368020 586168 368072 586220
rect 378232 586168 378284 586220
rect 388628 586168 388680 586220
rect 398840 586168 398892 586220
rect 409236 586168 409288 586220
rect 443000 586236 443052 586288
rect 456248 586372 456300 586424
rect 456340 586372 456392 586424
rect 463700 586440 463752 586492
rect 473912 586372 473964 586424
rect 476856 586372 476908 586424
rect 476948 586372 477000 586424
rect 485780 586440 485832 586492
rect 432788 586168 432840 586220
rect 292948 586100 293000 586152
rect 294328 586100 294380 586152
rect 533988 586100 534040 586152
rect 271144 586032 271196 586084
rect 509884 586032 509936 586084
rect 239956 585896 240008 585948
rect 250260 585896 250312 585948
rect 265992 585896 266044 585948
rect 313648 585964 313700 586016
rect 461676 585964 461728 586016
rect 288532 585896 288584 585948
rect 557908 585896 557960 585948
rect 318616 582904 318668 582956
rect 560852 582904 560904 582956
rect 26516 582360 26568 582412
rect 270040 582360 270092 582412
rect 27252 582292 27304 582344
rect 275928 582292 275980 582344
rect 24860 582224 24912 582276
rect 314292 582224 314344 582276
rect 319444 582224 319496 582276
rect 558460 582224 558512 582276
rect 275928 580660 275980 580712
rect 315028 580660 315080 580712
rect 24952 576988 25004 577040
rect 26516 577056 26568 577108
rect 317972 576240 318024 576292
rect 319444 576240 319496 576292
rect 317144 572636 317196 572688
rect 317972 572636 318024 572688
rect 270040 569576 270092 569628
rect 273812 569576 273864 569628
rect 273812 565836 273864 565888
rect 275284 565836 275336 565888
rect 275284 562776 275336 562828
rect 279608 562776 279660 562828
rect 315028 562300 315080 562352
rect 317144 562300 317196 562352
rect 309784 559308 309836 559360
rect 315028 559376 315080 559428
rect 279700 556452 279752 556504
rect 285496 556384 285548 556436
rect 285496 549720 285548 549772
rect 290648 549720 290700 549772
rect 269304 547612 269356 547664
rect 314200 547544 314252 547596
rect 318616 547544 318668 547596
rect 314292 544892 314344 544944
rect 315028 544892 315080 544944
rect 307668 544552 307720 544604
rect 309784 544552 309836 544604
rect 290648 540200 290700 540252
rect 293316 540132 293368 540184
rect 293316 537208 293368 537260
rect 294420 537208 294472 537260
rect 304724 536528 304776 536580
rect 307668 536528 307720 536580
rect 303252 534488 303304 534540
rect 304724 534488 304776 534540
rect 294420 534352 294472 534404
rect 298008 534216 298060 534268
rect 298836 529864 298888 529916
rect 303252 529932 303304 529984
rect 298008 523948 298060 524000
rect 300124 523948 300176 524000
rect 295064 522588 295116 522640
rect 298744 522588 298796 522640
rect 300124 519052 300176 519104
rect 301596 519052 301648 519104
rect 301596 516672 301648 516724
rect 303160 516672 303212 516724
rect 303160 515176 303212 515228
rect 307392 515108 307444 515160
rect 558460 512116 558512 512168
rect 558920 512116 558972 512168
rect 269304 511504 269356 511556
rect 272156 511504 272208 511556
rect 295064 511504 295116 511556
rect 307392 509668 307444 509720
rect 315028 509668 315080 509720
rect 307392 487228 307444 487280
rect 307576 487228 307628 487280
rect 2964 479884 3016 479936
rect 3976 479884 4028 479936
rect 270040 472540 270092 472592
rect 315028 472540 315080 472592
rect 307392 466624 307444 466676
rect 307576 466624 307628 466676
rect 307392 446020 307444 446072
rect 307576 446020 307628 446072
rect 558460 440444 558512 440496
rect 558920 440444 558972 440496
rect 269304 440104 269356 440156
rect 286232 440104 286284 440156
rect 307392 425416 307444 425468
rect 307576 425416 307628 425468
rect 269304 404812 269356 404864
rect 303896 404812 303948 404864
rect 298744 386384 298796 386436
rect 298836 386384 298888 386436
rect 24952 386180 25004 386232
rect 278136 386248 278188 386300
rect 291384 386316 291436 386368
rect 309048 386316 309100 386368
rect 314384 386316 314436 386368
rect 286232 386248 286284 386300
rect 558460 386248 558512 386300
rect 267924 386180 267976 386232
rect 291384 386112 291436 386164
rect 298744 386112 298796 386164
rect 314016 385704 314068 385756
rect 314384 385704 314436 385756
rect 303896 384888 303948 384940
rect 312636 384888 312688 384940
rect 560852 384888 560904 384940
rect 307392 384208 307444 384260
rect 307576 384208 307628 384260
rect 256056 382644 256108 382696
rect 271052 382644 271104 382696
rect 275284 382644 275336 382696
rect 286324 382644 286376 382696
rect 301688 382644 301740 382696
rect 331496 382644 331548 382696
rect 232136 382576 232188 382628
rect 313556 382576 313608 382628
rect 270132 382508 270184 382560
rect 355600 382508 355652 382560
rect 270960 382440 271012 382492
rect 271972 382440 272024 382492
rect 379520 382440 379572 382492
rect 208032 382372 208084 382424
rect 278228 382372 278280 382424
rect 279516 382372 279568 382424
rect 279700 382372 279752 382424
rect 403624 382372 403676 382424
rect 183928 382304 183980 382356
rect 264980 382304 265032 382356
rect 275192 382304 275244 382356
rect 275284 382304 275336 382356
rect 111800 382236 111852 382288
rect 279700 382236 279752 382288
rect 286324 382236 286376 382288
rect 295892 382236 295944 382288
rect 316408 382236 316460 382288
rect 475936 382236 475988 382288
rect 135904 382168 135956 382220
rect 314108 382168 314160 382220
rect 427728 382168 427780 382220
rect 87696 382100 87748 382152
rect 270960 382100 271012 382152
rect 279516 382100 279568 382152
rect 499856 382100 499908 382152
rect 39672 382032 39724 382084
rect 301688 382032 301740 382084
rect 313556 382032 313608 382084
rect 313924 382032 313976 382084
rect 523960 382032 524012 382084
rect 63776 381964 63828 382016
rect 270132 381964 270184 382016
rect 271052 381964 271104 382016
rect 272064 381964 272116 382016
rect 548064 381964 548116 382016
rect 264980 381896 265032 381948
rect 275192 381896 275244 381948
rect 295892 381896 295944 381948
rect 313832 381896 313884 381948
rect 316408 381896 316460 381948
rect 273168 359388 273220 359440
rect 278596 359388 278648 359440
rect 273352 359320 273404 359372
rect 286232 359320 286284 359372
rect 301228 359320 301280 359372
rect 301688 359320 301740 359372
rect 306932 359388 306984 359440
rect 307024 359388 307076 359440
rect 312544 359388 312596 359440
rect 306932 359252 306984 359304
rect 312268 359252 312320 359304
rect 273444 359184 273496 359236
rect 278504 359184 278556 359236
rect 278596 359184 278648 359236
rect 288808 359184 288860 359236
rect 292948 359184 293000 359236
rect 294328 359184 294380 359236
rect 307024 359184 307076 359236
rect 307576 359184 307628 359236
rect 312452 359184 312504 359236
rect 305276 358504 305328 358556
rect 579252 358504 579304 358556
rect 267096 358436 267148 358488
rect 294972 358436 295024 358488
rect 303252 358436 303304 358488
rect 579344 358436 579396 358488
rect 3976 358368 4028 358420
rect 274364 358368 274416 358420
rect 282644 358368 282696 358420
rect 579620 358368 579672 358420
rect 299020 358300 299072 358352
rect 300216 358300 300268 358352
rect 24952 357892 25004 357944
rect 311348 357892 311400 357944
rect 271512 357824 271564 357876
rect 296996 357824 297048 357876
rect 147128 357756 147180 357808
rect 284668 357756 284720 357808
rect 290924 357756 290976 357808
rect 317144 357756 317196 357808
rect 309324 357688 309376 357740
rect 315672 357688 315724 357740
rect 273260 356260 273312 356312
rect 275928 356260 275980 356312
rect 273536 354832 273588 354884
rect 279700 354832 279752 354884
rect 280252 354832 280304 354884
rect 3884 354084 3936 354136
rect 311532 354084 311584 354136
rect 270316 354016 270368 354068
rect 579436 354016 579488 354068
rect 3792 353948 3844 354000
rect 313556 353948 313608 354000
rect 269856 353200 269908 353252
rect 270132 353200 270184 353252
rect 269672 350276 269724 350328
rect 269856 350276 269908 350328
rect 269672 340076 269724 340128
rect 269948 340008 270000 340060
rect 268568 339940 268620 339992
rect 269672 339940 269724 339992
rect 314016 334092 314068 334144
rect 579160 334092 579212 334144
rect 314016 333412 314068 333464
rect 314292 333412 314344 333464
rect 268568 329740 268620 329792
rect 269396 329740 269448 329792
rect 272156 316208 272208 316260
rect 275284 316208 275336 316260
rect 310888 316208 310940 316260
rect 312728 316208 312780 316260
rect 3608 313488 3660 313540
rect 308588 313488 308640 313540
rect 3700 313420 3752 313472
rect 285956 313420 286008 313472
rect 287980 313420 288032 313472
rect 579528 313420 579580 313472
rect 272248 313352 272300 313404
rect 283932 313352 283984 313404
rect 292212 313352 292264 313404
rect 561496 313352 561548 313404
rect 24860 313284 24912 313336
rect 273628 313284 273680 313336
rect 277676 313284 277728 313336
rect 312820 313284 312872 313336
rect 271972 313216 272024 313268
rect 281908 313216 281960 313268
rect 296260 313216 296312 313268
rect 297272 313216 297324 313268
rect 313924 313216 313976 313268
rect 272064 313148 272116 313200
rect 279700 313148 279752 313200
rect 298744 313148 298796 313200
rect 313648 313148 313700 313200
rect 306564 313012 306616 313064
rect 307576 313012 307628 313064
rect 313740 313012 313792 313064
rect 122104 312876 122156 312928
rect 290004 312876 290056 312928
rect 98552 312808 98604 312860
rect 300308 312808 300360 312860
rect 24860 312740 24912 312792
rect 302516 312740 302568 312792
rect 270040 312128 270092 312180
rect 281172 312060 281224 312112
rect 281908 312060 281960 312112
rect 282644 312060 282696 312112
rect 283932 312060 283984 312112
rect 270040 311992 270092 312044
rect 303896 311992 303948 312044
rect 304540 311992 304592 312044
rect 312636 311992 312688 312044
rect 270040 309068 270092 309120
rect 270316 309068 270368 309120
rect 269856 291456 269908 291508
rect 269948 291320 270000 291372
rect 98000 276700 98052 276752
rect 98552 276700 98604 276752
rect 146208 276700 146260 276752
rect 147128 276700 147180 276752
rect 170128 276632 170180 276684
rect 175188 276632 175240 276684
rect 185400 276564 185452 276616
rect 188344 276564 188396 276616
rect 188436 276564 188488 276616
rect 195796 276632 195848 276684
rect 206008 276564 206060 276616
rect 208952 276564 209004 276616
rect 209044 276564 209096 276616
rect 216404 276632 216456 276684
rect 226616 276564 226668 276616
rect 229560 276564 229612 276616
rect 229652 276564 229704 276616
rect 237012 276632 237064 276684
rect 257620 276632 257672 276684
rect 267832 276632 267884 276684
rect 240048 276564 240100 276616
rect 250260 276564 250312 276616
rect 285588 276564 285640 276616
rect 295800 276564 295852 276616
rect 307024 276564 307076 276616
rect 307576 276564 307628 276616
rect 341800 276564 341852 276616
rect 242440 276496 242492 276548
rect 312084 276496 312136 276548
rect 312544 276496 312596 276548
rect 326896 276496 326948 276548
rect 337016 276496 337068 276548
rect 347504 276496 347556 276548
rect 357624 276496 357676 276548
rect 257620 276428 257672 276480
rect 267832 276428 267884 276480
rect 250260 276360 250312 276412
rect 282644 276428 282696 276480
rect 365720 276496 365772 276548
rect 403992 276496 404044 276548
rect 419448 276496 419500 276548
rect 362776 276428 362828 276480
rect 378232 276428 378284 276480
rect 383384 276428 383436 276480
rect 398840 276428 398892 276480
rect 429844 276428 429896 276480
rect 435640 276428 435692 276480
rect 435732 276428 435784 276480
rect 443092 276496 443144 276548
rect 453304 276428 453356 276480
rect 454224 276428 454276 276480
rect 294328 276360 294380 276412
rect 413928 276360 413980 276412
rect 285588 276292 285640 276344
rect 317144 276292 317196 276344
rect 438032 276292 438084 276344
rect 73528 276224 73580 276276
rect 282644 276224 282696 276276
rect 295800 276224 295852 276276
rect 298744 276224 298796 276276
rect 306196 276224 306248 276276
rect 316408 276224 316460 276276
rect 326896 276224 326948 276276
rect 337016 276224 337068 276276
rect 347504 276224 347556 276276
rect 357624 276224 357676 276276
rect 362776 276224 362828 276276
rect 378232 276224 378284 276276
rect 383384 276224 383436 276276
rect 398840 276224 398892 276276
rect 403992 276224 404044 276276
rect 419448 276224 419500 276276
rect 429844 276224 429896 276276
rect 454224 276224 454276 276276
rect 461952 276224 462004 276276
rect 194232 276156 194284 276208
rect 270408 276156 270460 276208
rect 486056 276156 486108 276208
rect 218336 276088 218388 276140
rect 270224 276088 270276 276140
rect 510160 276088 510212 276140
rect 49976 276020 50028 276072
rect 307024 276020 307076 276072
rect 312084 276020 312136 276072
rect 534264 276020 534316 276072
rect 266360 275952 266412 276004
rect 273168 275952 273220 276004
rect 558184 275952 558236 276004
rect 306196 275884 306248 275936
rect 316408 275884 316460 275936
rect 314384 272348 314436 272400
rect 560852 272348 560904 272400
rect 275928 272212 275980 272264
rect 26424 272076 26476 272128
rect 273260 272076 273312 272128
rect 276664 272076 276716 272128
rect 558644 272076 558696 272128
rect 27160 272008 27212 272060
rect 312544 272008 312596 272060
rect 27620 271940 27672 271992
rect 314016 271940 314068 271992
rect 314016 270852 314068 270904
rect 314292 270852 314344 270904
rect 276664 270784 276716 270836
rect 315028 270784 315080 270836
rect 26148 267928 26200 267980
rect 27620 267928 27672 267980
rect 558460 267928 558512 267980
rect 558644 267928 558696 267980
rect 558552 257524 558604 257576
rect 558644 257524 558696 257576
rect 24768 256164 24820 256216
rect 27160 256164 27212 256216
rect 558552 247256 558604 247308
rect 558736 247256 558788 247308
rect 268384 238416 268436 238468
rect 314384 238416 314436 238468
rect 270132 236988 270184 237040
rect 270224 236988 270276 237040
rect 558552 236988 558604 237040
rect 558828 236988 558880 237040
rect 558828 229712 558880 229764
rect 558736 229576 558788 229628
rect 269856 226720 269908 226772
rect 270224 226720 270276 226772
rect 270132 216384 270184 216436
rect 270224 216384 270276 216436
rect 270224 206048 270276 206100
rect 270408 206048 270460 206100
rect 558460 203124 558512 203176
rect 558828 203124 558880 203176
rect 268384 202784 268436 202836
rect 275928 202784 275980 202836
rect 312728 200132 312780 200184
rect 315028 200132 315080 200184
rect 270132 195780 270184 195832
rect 270408 195780 270460 195832
rect 270224 185444 270276 185496
rect 270408 185444 270460 185496
rect 270132 175176 270184 175228
rect 270408 175176 270460 175228
rect 270224 164772 270276 164824
rect 270408 164772 270460 164824
rect 270132 147296 270184 147348
rect 270132 147160 270184 147212
rect 270132 144236 270184 144288
rect 270224 144236 270276 144288
rect 270132 142740 270184 142792
rect 270408 142740 270460 142792
rect 270132 132472 270184 132524
rect 270224 132404 270276 132456
rect 268292 130568 268344 130620
rect 273352 130568 273404 130620
rect 273352 130228 273404 130280
rect 291476 130228 291528 130280
rect 270132 126624 270184 126676
rect 270224 126488 270276 126540
rect 558552 125604 558604 125656
rect 559380 125604 559432 125656
rect 291476 125536 291528 125588
rect 293592 125536 293644 125588
rect 270224 116288 270276 116340
rect 293592 116220 293644 116272
rect 294696 116220 294748 116272
rect 270316 116152 270368 116204
rect 294696 114724 294748 114776
rect 296444 114724 296496 114776
rect 296444 111800 296496 111852
rect 297364 111800 297416 111852
rect 297364 109284 297416 109336
rect 300216 109284 300268 109336
rect 270224 101600 270276 101652
rect 270316 101600 270368 101652
rect 300308 101532 300360 101584
rect 301780 101532 301832 101584
rect 267924 94868 267976 94920
rect 303896 94868 303948 94920
rect 301780 94188 301832 94240
rect 304724 94120 304776 94172
rect 314200 92352 314252 92404
rect 315028 92352 315080 92404
rect 269948 91264 270000 91316
rect 270132 91264 270184 91316
rect 304724 90380 304776 90432
rect 307668 90380 307720 90432
rect 307668 86844 307720 86896
rect 312084 86776 312136 86828
rect 269948 82424 270000 82476
rect 270316 82424 270368 82476
rect 312084 81132 312136 81184
rect 316500 81132 316552 81184
rect 24952 75964 25004 76016
rect 314200 75964 314252 76016
rect 316500 75964 316552 76016
rect 558552 75964 558604 76016
rect 303896 75896 303948 75948
rect 560852 75896 560904 75948
rect 39672 72088 39724 72140
rect 312360 72088 312412 72140
rect 313556 72088 313608 72140
rect 475936 72088 475988 72140
rect 63776 72020 63828 72072
rect 269396 72020 269448 72072
rect 279700 72020 279752 72072
rect 280160 72020 280212 72072
rect 548064 72020 548116 72072
rect 272340 71952 272392 72004
rect 273444 71952 273496 72004
rect 499856 71952 499908 72004
rect 87696 71884 87748 71936
rect 281172 71884 281224 71936
rect 297272 71884 297324 71936
rect 523960 71884 524012 71936
rect 135904 71816 135956 71868
rect 314108 71816 314160 71868
rect 427728 71816 427780 71868
rect 183928 71748 183980 71800
rect 313556 71748 313608 71800
rect 160008 71680 160060 71732
rect 271512 71680 271564 71732
rect 272432 71680 272484 71732
rect 273536 71680 273588 71732
rect 403624 71680 403676 71732
rect 208032 71612 208084 71664
rect 272340 71612 272392 71664
rect 281172 71612 281224 71664
rect 379520 71612 379572 71664
rect 269396 71544 269448 71596
rect 270316 71544 270368 71596
rect 355600 71544 355652 71596
rect 232136 71476 232188 71528
rect 297272 71476 297324 71528
rect 312360 71476 312412 71528
rect 331496 71476 331548 71528
rect 256056 71408 256108 71460
rect 280160 71408 280212 71460
rect 111800 71340 111852 71392
rect 272432 71340 272484 71392
rect 270592 3612 270644 3664
rect 583392 3612 583444 3664
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 703474 8156 703520
rect 8128 703446 8248 703474
rect 8220 700670 8248 703446
rect 8024 700664 8076 700670
rect 8024 700606 8076 700612
rect 8208 700664 8260 700670
rect 8208 700606 8260 700612
rect 3606 667992 3662 668001
rect 3606 667927 3662 667936
rect 2962 653576 3018 653585
rect 2962 653511 2964 653520
rect 3016 653511 3018 653520
rect 2964 653482 3016 653488
rect 2976 596057 3004 653482
rect 2962 596048 3018 596057
rect 2962 595983 3018 595992
rect 2976 538665 3004 595983
rect 2962 538656 3018 538665
rect 2962 538591 3018 538600
rect 2976 481137 3004 538591
rect 2962 481128 3018 481137
rect 2962 481063 3018 481072
rect 2976 479942 3004 481063
rect 2964 479936 3016 479942
rect 2964 479878 3016 479884
rect 3620 313546 3648 667927
rect 8036 653546 8064 700606
rect 24320 699922 24348 703520
rect 72988 700670 73016 703520
rect 72976 700664 73028 700670
rect 72976 700606 73028 700612
rect 89180 700058 89208 703520
rect 137848 700670 137876 703520
rect 137836 700664 137888 700670
rect 137836 700606 137888 700612
rect 89168 700052 89220 700058
rect 89168 699994 89220 700000
rect 154132 699990 154160 703520
rect 202800 700670 202828 703520
rect 202788 700664 202840 700670
rect 202788 700606 202840 700612
rect 218992 700194 219020 703520
rect 267660 700670 267688 703520
rect 267648 700664 267700 700670
rect 267648 700606 267700 700612
rect 283852 700330 283880 703520
rect 332520 700670 332548 703520
rect 332508 700664 332560 700670
rect 332508 700606 332560 700612
rect 272984 700324 273036 700330
rect 272984 700266 273036 700272
rect 283840 700324 283892 700330
rect 283840 700266 283892 700272
rect 270868 700256 270920 700262
rect 270868 700198 270920 700204
rect 218980 700188 219032 700194
rect 218980 700130 219032 700136
rect 270684 700120 270736 700126
rect 270684 700062 270736 700068
rect 154120 699984 154172 699990
rect 154120 699926 154172 699932
rect 268568 699984 268620 699990
rect 268568 699926 268620 699932
rect 24308 699916 24360 699922
rect 24308 699858 24360 699864
rect 8024 653540 8076 653546
rect 8024 653482 8076 653488
rect 3698 610464 3754 610473
rect 3698 610399 3754 610408
rect 3608 313540 3660 313546
rect 3608 313482 3660 313488
rect 3712 313478 3740 610399
rect 49608 586628 49660 586634
rect 49608 586570 49660 586576
rect 49620 583930 49648 586570
rect 217968 586560 218020 586566
rect 217968 586502 218020 586508
rect 73528 586492 73580 586498
rect 73528 586434 73580 586440
rect 73540 583930 73568 586434
rect 169760 586356 169812 586362
rect 169760 586298 169812 586304
rect 121736 586288 121788 586294
rect 121736 586230 121788 586236
rect 121748 583930 121776 586230
rect 145840 586084 145892 586090
rect 145840 586026 145892 586032
rect 145852 583930 145880 586026
rect 169772 583930 169800 586298
rect 198740 586220 198792 586226
rect 198740 586162 198792 586168
rect 209044 586220 209096 586226
rect 209044 586162 209096 586168
rect 216496 586220 216548 586226
rect 216496 586162 216548 586168
rect 198752 586022 198780 586162
rect 193864 586016 193916 586022
rect 193864 585958 193916 585964
rect 198740 586016 198792 586022
rect 198740 585958 198792 585964
rect 193876 583930 193904 585958
rect 209056 585954 209084 586162
rect 209044 585948 209096 585954
rect 209044 585890 209096 585896
rect 216404 585948 216456 585954
rect 216404 585890 216456 585896
rect 216416 585834 216444 585890
rect 216508 585834 216536 586162
rect 216416 585806 216536 585834
rect 217980 583930 218008 586502
rect 242072 586424 242124 586430
rect 242072 586366 242124 586372
rect 229652 586220 229704 586226
rect 229652 586162 229704 586168
rect 229664 586022 229692 586162
rect 239956 586152 240008 586158
rect 239956 586094 240008 586100
rect 229652 586016 229704 586022
rect 229652 585958 229704 585964
rect 239968 585954 239996 586094
rect 239956 585948 240008 585954
rect 239956 585890 240008 585896
rect 242084 583930 242112 586366
rect 250260 586152 250312 586158
rect 250260 586094 250312 586100
rect 257618 586120 257674 586129
rect 250272 585954 250300 586094
rect 267738 586120 267794 586129
rect 257618 586055 257674 586064
rect 267096 586084 267148 586090
rect 257632 586022 257660 586055
rect 267738 586055 267794 586064
rect 267096 586026 267148 586032
rect 257620 586016 257672 586022
rect 257620 585958 257672 585964
rect 250260 585948 250312 585954
rect 250260 585890 250312 585896
rect 265992 585948 266044 585954
rect 265992 585890 266044 585896
rect 266004 583930 266032 585890
rect 49620 583902 49680 583930
rect 73540 583902 73600 583930
rect 121748 583902 121808 583930
rect 145852 583902 145912 583930
rect 169772 583902 169832 583930
rect 193876 583902 193936 583930
rect 217980 583902 218040 583930
rect 242084 583902 242144 583930
rect 266004 583902 266064 583930
rect 26516 582412 26568 582418
rect 26516 582354 26568 582360
rect 24860 582276 24912 582282
rect 24860 582218 24912 582224
rect 3790 553072 3846 553081
rect 3790 553007 3846 553016
rect 3804 354006 3832 553007
rect 24872 545601 24900 582218
rect 26528 577114 26556 582354
rect 27252 582344 27304 582350
rect 27252 582286 27304 582292
rect 27264 581233 27292 582286
rect 27250 581224 27306 581233
rect 27250 581159 27306 581168
rect 26516 577108 26568 577114
rect 26516 577050 26568 577056
rect 24952 577040 25004 577046
rect 24952 576982 25004 576988
rect 24858 545592 24914 545601
rect 24858 545527 24914 545536
rect 24964 509969 24992 576982
rect 24950 509960 25006 509969
rect 24950 509895 25006 509904
rect 3882 495544 3938 495553
rect 3882 495479 3938 495488
rect 3896 354142 3924 495479
rect 3976 479936 4028 479942
rect 3976 479878 4028 479884
rect 3988 358426 4016 479878
rect 24858 473104 24914 473113
rect 24858 473039 24914 473048
rect 3976 358420 4028 358426
rect 3976 358362 4028 358368
rect 3884 354136 3936 354142
rect 3884 354078 3936 354084
rect 3792 354000 3844 354006
rect 3792 353942 3844 353948
rect 3700 313472 3752 313478
rect 3700 313414 3752 313420
rect 24872 313342 24900 473039
rect 24950 402112 25006 402121
rect 24950 402047 25006 402056
rect 24964 386238 24992 402047
rect 24952 386232 25004 386238
rect 24952 386174 25004 386180
rect 39376 383982 39712 384010
rect 63480 383982 63816 384010
rect 87400 383982 87736 384010
rect 111504 383982 111840 384010
rect 135608 383982 135944 384010
rect 183816 383982 183968 384010
rect 207736 383982 208072 384010
rect 231840 383982 232176 384010
rect 255944 383982 256096 384010
rect 39684 382090 39712 383982
rect 39672 382084 39724 382090
rect 39672 382026 39724 382032
rect 63788 382022 63816 383982
rect 87708 382158 87736 383982
rect 111812 382294 111840 383982
rect 111800 382288 111852 382294
rect 111800 382230 111852 382236
rect 135916 382226 135944 383982
rect 183940 382362 183968 383982
rect 208044 382430 208072 383982
rect 232148 382634 232176 383982
rect 256068 382702 256096 383982
rect 256056 382696 256108 382702
rect 256056 382638 256108 382644
rect 232136 382628 232188 382634
rect 232136 382570 232188 382576
rect 208032 382424 208084 382430
rect 208032 382366 208084 382372
rect 183928 382356 183980 382362
rect 183928 382298 183980 382304
rect 264980 382356 265032 382362
rect 264980 382298 265032 382304
rect 135904 382220 135956 382226
rect 135904 382162 135956 382168
rect 87696 382152 87748 382158
rect 87696 382094 87748 382100
rect 63776 382016 63828 382022
rect 63776 381958 63828 381964
rect 264992 381954 265020 382298
rect 264980 381948 265032 381954
rect 264980 381890 265032 381896
rect 267108 358494 267136 586026
rect 267752 586022 267780 586055
rect 267740 586016 267792 586022
rect 267740 585958 267792 585964
rect 267924 386232 267976 386238
rect 267922 386200 267924 386209
rect 267976 386200 267978 386209
rect 267922 386135 267978 386144
rect 267096 358488 267148 358494
rect 267096 358430 267148 358436
rect 24952 357944 25004 357950
rect 24952 357886 25004 357892
rect 24860 313336 24912 313342
rect 24860 313278 24912 313284
rect 24860 312792 24912 312798
rect 24860 312734 24912 312740
rect 24768 256216 24820 256222
rect 24768 256158 24820 256164
rect 24780 199073 24808 256158
rect 24766 199064 24822 199073
rect 24766 198999 24822 199008
rect 24872 163441 24900 312734
rect 24858 163432 24914 163441
rect 24858 163367 24914 163376
rect 24964 128081 24992 357886
rect 147128 357808 147180 357814
rect 147128 357750 147180 357756
rect 122104 312928 122156 312934
rect 122104 312870 122156 312876
rect 98552 312860 98604 312866
rect 98552 312802 98604 312808
rect 98564 276758 98592 312802
rect 98000 276752 98052 276758
rect 98000 276694 98052 276700
rect 98552 276752 98604 276758
rect 98552 276694 98604 276700
rect 73528 276276 73580 276282
rect 73528 276218 73580 276224
rect 49976 276072 50028 276078
rect 49976 276014 50028 276020
rect 49988 273578 50016 276014
rect 49680 273550 50016 273578
rect 73540 273578 73568 276218
rect 98012 273578 98040 276694
rect 122116 273578 122144 312870
rect 147140 276758 147168 357750
rect 268580 339998 268608 699926
rect 270500 627156 270552 627162
rect 270500 627098 270552 627104
rect 270408 586152 270460 586158
rect 270408 586094 270460 586100
rect 270040 582412 270092 582418
rect 270040 582354 270092 582360
rect 270052 569634 270080 582354
rect 270040 569628 270092 569634
rect 270040 569570 270092 569576
rect 269304 547664 269356 547670
rect 269302 547632 269304 547641
rect 269356 547632 269358 547641
rect 269302 547567 269358 547576
rect 269302 512000 269358 512009
rect 269302 511935 269358 511944
rect 269316 511562 269344 511935
rect 269304 511556 269356 511562
rect 269304 511498 269356 511504
rect 270040 472592 270092 472598
rect 270040 472534 270092 472540
rect 269302 440736 269358 440745
rect 269302 440671 269358 440680
rect 269316 440162 269344 440671
rect 269304 440156 269356 440162
rect 269304 440098 269356 440104
rect 269302 405376 269358 405385
rect 269302 405311 269358 405320
rect 269316 404870 269344 405311
rect 269304 404864 269356 404870
rect 269304 404806 269356 404812
rect 269856 353252 269908 353258
rect 269856 353194 269908 353200
rect 269868 350334 269896 353194
rect 269672 350328 269724 350334
rect 269672 350270 269724 350276
rect 269856 350328 269908 350334
rect 269856 350270 269908 350276
rect 269684 340134 269712 350270
rect 270052 348809 270080 472534
rect 270132 382560 270184 382566
rect 270132 382502 270184 382508
rect 270144 382022 270172 382502
rect 270132 382016 270184 382022
rect 270132 381958 270184 381964
rect 270144 353258 270172 381958
rect 270316 354068 270368 354074
rect 270316 354010 270368 354016
rect 270222 353832 270278 353841
rect 270222 353767 270278 353776
rect 270132 353252 270184 353258
rect 270132 353194 270184 353200
rect 270038 348800 270094 348809
rect 270038 348735 270094 348744
rect 269672 340128 269724 340134
rect 269672 340070 269724 340076
rect 269948 340060 270000 340066
rect 269948 340002 270000 340008
rect 268568 339992 268620 339998
rect 268568 339934 268620 339940
rect 269672 339992 269724 339998
rect 269960 339969 269988 340002
rect 269672 339934 269724 339940
rect 269946 339960 270002 339969
rect 269684 339697 269712 339934
rect 269946 339895 270002 339904
rect 270130 339824 270186 339833
rect 270130 339759 270186 339768
rect 269670 339688 269726 339697
rect 269670 339623 269726 339632
rect 270144 335617 270172 339759
rect 269854 335608 269910 335617
rect 269854 335543 269910 335552
rect 270130 335608 270186 335617
rect 270130 335543 270186 335552
rect 269394 329896 269450 329905
rect 269394 329831 269450 329840
rect 269408 329798 269436 329831
rect 268568 329792 268620 329798
rect 268568 329734 268620 329740
rect 269396 329792 269448 329798
rect 269396 329734 269448 329740
rect 146208 276752 146260 276758
rect 146208 276694 146260 276700
rect 147128 276752 147180 276758
rect 147128 276694 147180 276700
rect 175186 276720 175242 276729
rect 146220 273578 146248 276694
rect 170128 276684 170180 276690
rect 175186 276655 175188 276664
rect 170128 276626 170180 276632
rect 175240 276655 175242 276664
rect 185398 276720 185454 276729
rect 185398 276655 185454 276664
rect 195794 276720 195850 276729
rect 195794 276655 195796 276664
rect 175188 276626 175240 276632
rect 170140 273578 170168 276626
rect 185412 276622 185440 276655
rect 195848 276655 195850 276664
rect 206006 276720 206062 276729
rect 206006 276655 206062 276664
rect 216402 276720 216458 276729
rect 216402 276655 216404 276664
rect 195796 276626 195848 276632
rect 206020 276622 206048 276655
rect 216456 276655 216458 276664
rect 226614 276720 226670 276729
rect 226614 276655 226670 276664
rect 237010 276720 237066 276729
rect 237010 276655 237012 276664
rect 216404 276626 216456 276632
rect 226628 276622 226656 276655
rect 237064 276655 237066 276664
rect 240046 276720 240102 276729
rect 240046 276655 240102 276664
rect 257620 276684 257672 276690
rect 237012 276626 237064 276632
rect 240060 276622 240088 276655
rect 257620 276626 257672 276632
rect 267832 276684 267884 276690
rect 267832 276626 267884 276632
rect 185400 276616 185452 276622
rect 185400 276558 185452 276564
rect 188344 276616 188396 276622
rect 188436 276616 188488 276622
rect 188396 276564 188436 276570
rect 188344 276558 188488 276564
rect 206008 276616 206060 276622
rect 206008 276558 206060 276564
rect 208952 276616 209004 276622
rect 209044 276616 209096 276622
rect 209004 276564 209044 276570
rect 208952 276558 209096 276564
rect 226616 276616 226668 276622
rect 226616 276558 226668 276564
rect 229560 276616 229612 276622
rect 229652 276616 229704 276622
rect 229612 276564 229652 276570
rect 229560 276558 229704 276564
rect 240048 276616 240100 276622
rect 240048 276558 240100 276564
rect 250260 276616 250312 276622
rect 250260 276558 250312 276564
rect 188356 276542 188476 276558
rect 208964 276542 209084 276558
rect 229572 276542 229692 276558
rect 242440 276548 242492 276554
rect 242440 276490 242492 276496
rect 194232 276208 194284 276214
rect 194232 276150 194284 276156
rect 194244 273578 194272 276150
rect 218336 276140 218388 276146
rect 218336 276082 218388 276088
rect 218348 273578 218376 276082
rect 242452 273578 242480 276490
rect 250272 276418 250300 276558
rect 257632 276486 257660 276626
rect 267844 276486 267872 276626
rect 257620 276480 257672 276486
rect 257620 276422 257672 276428
rect 267832 276480 267884 276486
rect 267832 276422 267884 276428
rect 250260 276412 250312 276418
rect 250260 276354 250312 276360
rect 266360 276004 266412 276010
rect 266360 275946 266412 275952
rect 266372 273578 266400 275946
rect 73540 273550 73600 273578
rect 97704 273550 98040 273578
rect 121808 273550 122144 273578
rect 145912 273550 146248 273578
rect 169832 273550 170168 273578
rect 193936 273550 194272 273578
rect 218040 273550 218376 273578
rect 242144 273550 242480 273578
rect 266064 273550 266400 273578
rect 26424 272128 26476 272134
rect 26424 272070 26476 272076
rect 26436 270337 26464 272070
rect 27160 272060 27212 272066
rect 27160 272002 27212 272008
rect 26422 270328 26478 270337
rect 26422 270263 26478 270272
rect 26148 267980 26200 267986
rect 26148 267922 26200 267928
rect 26160 260522 26188 267922
rect 26160 260494 26280 260522
rect 26252 250322 26280 260494
rect 27172 256222 27200 272002
rect 27620 271992 27672 271998
rect 27620 271934 27672 271940
rect 27632 267986 27660 271934
rect 27620 267980 27672 267986
rect 27620 267922 27672 267928
rect 27160 256216 27212 256222
rect 27160 256158 27212 256164
rect 26252 250294 26372 250322
rect 26344 239986 26372 250294
rect 26344 239958 26464 239986
rect 26436 234705 26464 239958
rect 268384 238468 268436 238474
rect 268384 238410 268436 238416
rect 268396 237425 268424 238410
rect 268382 237416 268438 237425
rect 268382 237351 268438 237360
rect 26422 234696 26478 234705
rect 26422 234631 26478 234640
rect 268384 202836 268436 202842
rect 268384 202778 268436 202784
rect 268396 201793 268424 202778
rect 268382 201784 268438 201793
rect 268382 201719 268438 201728
rect 268580 166161 268608 329734
rect 269868 322402 269896 335543
rect 269868 322374 270080 322402
rect 270052 312186 270080 322374
rect 270040 312180 270092 312186
rect 270040 312122 270092 312128
rect 270040 312044 270092 312050
rect 270040 311986 270092 311992
rect 270052 309126 270080 311986
rect 270040 309120 270092 309126
rect 270040 309062 270092 309068
rect 269854 297392 269910 297401
rect 269854 297327 269910 297336
rect 269868 291514 269896 297327
rect 269856 291508 269908 291514
rect 269856 291450 269908 291456
rect 269948 291372 270000 291378
rect 269948 291314 270000 291320
rect 269960 260522 269988 291314
rect 270236 276146 270264 353767
rect 270328 324465 270356 354010
rect 270420 345273 270448 586094
rect 270406 345264 270462 345273
rect 270406 345199 270462 345208
rect 270314 324456 270370 324465
rect 270314 324391 270370 324400
rect 270316 309120 270368 309126
rect 270316 309062 270368 309068
rect 270328 297401 270356 309062
rect 270314 297392 270370 297401
rect 270314 297327 270370 297336
rect 270420 276214 270448 345199
rect 270512 320793 270540 627098
rect 270592 586560 270644 586566
rect 270592 586502 270644 586508
rect 270604 353841 270632 586502
rect 270590 353832 270646 353841
rect 270590 353767 270646 353776
rect 270590 350840 270646 350849
rect 270590 350775 270646 350784
rect 270498 320784 270554 320793
rect 270498 320719 270554 320728
rect 270408 276208 270460 276214
rect 270408 276150 270460 276156
rect 270224 276140 270276 276146
rect 270224 276082 270276 276088
rect 269960 260494 270080 260522
rect 270052 250322 270080 260494
rect 270052 250294 270264 250322
rect 270144 237046 270172 237077
rect 270236 237046 270264 250294
rect 270132 237040 270184 237046
rect 269854 237008 269910 237017
rect 269854 236943 269910 236952
rect 270038 237008 270094 237017
rect 270094 236988 270132 236994
rect 270094 236982 270184 236988
rect 270224 237040 270276 237046
rect 270224 236982 270276 236988
rect 270094 236966 270172 236982
rect 270038 236943 270094 236952
rect 269868 226778 269896 236943
rect 269856 226772 269908 226778
rect 269856 226714 269908 226720
rect 270224 226772 270276 226778
rect 270224 226714 270276 226720
rect 270236 216442 270264 226714
rect 270132 216436 270184 216442
rect 270132 216378 270184 216384
rect 270224 216436 270276 216442
rect 270224 216378 270276 216384
rect 270144 209114 270172 216378
rect 270144 209086 270264 209114
rect 270236 206106 270264 209086
rect 270224 206100 270276 206106
rect 270224 206042 270276 206048
rect 270408 206100 270460 206106
rect 270408 206042 270460 206048
rect 270420 195838 270448 206042
rect 270132 195832 270184 195838
rect 270132 195774 270184 195780
rect 270408 195832 270460 195838
rect 270408 195774 270460 195780
rect 270144 188442 270172 195774
rect 270144 188414 270264 188442
rect 270236 185502 270264 188414
rect 270224 185496 270276 185502
rect 270224 185438 270276 185444
rect 270408 185496 270460 185502
rect 270408 185438 270460 185444
rect 270420 175234 270448 185438
rect 270132 175228 270184 175234
rect 270132 175170 270184 175176
rect 270408 175228 270460 175234
rect 270408 175170 270460 175176
rect 270144 167906 270172 175170
rect 270144 167878 270264 167906
rect 268566 166152 268622 166161
rect 268566 166087 268622 166096
rect 270236 164830 270264 167878
rect 270224 164824 270276 164830
rect 270224 164766 270276 164772
rect 270408 164824 270460 164830
rect 270408 164766 270460 164772
rect 270420 154601 270448 164766
rect 270130 154592 270186 154601
rect 270130 154527 270186 154536
rect 270406 154592 270462 154601
rect 270406 154527 270462 154536
rect 270144 147354 270172 154527
rect 270132 147348 270184 147354
rect 270132 147290 270184 147296
rect 270132 147212 270184 147218
rect 270132 147154 270184 147160
rect 270144 144294 270172 147154
rect 270132 144288 270184 144294
rect 270224 144288 270276 144294
rect 270132 144230 270184 144236
rect 270222 144256 270224 144265
rect 270276 144256 270278 144265
rect 270222 144191 270278 144200
rect 270406 144256 270462 144265
rect 270406 144191 270462 144200
rect 270420 142798 270448 144191
rect 270132 142792 270184 142798
rect 270132 142734 270184 142740
rect 270408 142792 270460 142798
rect 270408 142734 270460 142740
rect 270144 132530 270172 142734
rect 270132 132524 270184 132530
rect 270132 132466 270184 132472
rect 270224 132456 270276 132462
rect 270224 132398 270276 132404
rect 270236 131050 270264 132398
rect 270144 131022 270264 131050
rect 268292 130620 268344 130626
rect 268292 130562 268344 130568
rect 268304 130529 268332 130562
rect 268290 130520 268346 130529
rect 268290 130455 268346 130464
rect 24950 128072 25006 128081
rect 24950 128007 25006 128016
rect 270144 126682 270172 131022
rect 270132 126676 270184 126682
rect 270132 126618 270184 126624
rect 270224 126540 270276 126546
rect 270224 126482 270276 126488
rect 270236 116346 270264 126482
rect 270224 116340 270276 116346
rect 270224 116282 270276 116288
rect 270316 116204 270368 116210
rect 270316 116146 270368 116152
rect 270328 101658 270356 116146
rect 270224 101652 270276 101658
rect 270224 101594 270276 101600
rect 270316 101652 270368 101658
rect 270316 101594 270368 101600
rect 270236 101538 270264 101594
rect 270144 101510 270264 101538
rect 267922 95160 267978 95169
rect 267922 95095 267978 95104
rect 267936 94926 267964 95095
rect 267924 94920 267976 94926
rect 267924 94862 267976 94868
rect 24950 92440 25006 92449
rect 24950 92375 25006 92384
rect 24964 76022 24992 92375
rect 270144 91322 270172 101510
rect 269948 91316 270000 91322
rect 269948 91258 270000 91264
rect 270132 91316 270184 91322
rect 270132 91258 270184 91264
rect 269960 82482 269988 91258
rect 269948 82476 270000 82482
rect 269948 82418 270000 82424
rect 270316 82476 270368 82482
rect 270316 82418 270368 82424
rect 24952 76016 25004 76022
rect 24952 75958 25004 75964
rect 39376 73630 39712 73658
rect 63480 73630 63816 73658
rect 87400 73630 87736 73658
rect 111504 73630 111840 73658
rect 135608 73630 135944 73658
rect 159712 73630 160048 73658
rect 183816 73630 183968 73658
rect 207736 73630 208072 73658
rect 231840 73630 232176 73658
rect 255944 73630 256096 73658
rect 39684 72146 39712 73630
rect 39672 72140 39724 72146
rect 39672 72082 39724 72088
rect 63788 72078 63816 73630
rect 63776 72072 63828 72078
rect 63776 72014 63828 72020
rect 87708 71942 87736 73630
rect 87696 71936 87748 71942
rect 87696 71878 87748 71884
rect 111812 71398 111840 73630
rect 135916 71874 135944 73630
rect 135904 71868 135956 71874
rect 135904 71810 135956 71816
rect 160020 71738 160048 73630
rect 183940 71806 183968 73630
rect 183928 71800 183980 71806
rect 183928 71742 183980 71748
rect 160008 71732 160060 71738
rect 160008 71674 160060 71680
rect 208044 71670 208072 73630
rect 208032 71664 208084 71670
rect 208032 71606 208084 71612
rect 232148 71534 232176 73630
rect 232136 71528 232188 71534
rect 232136 71470 232188 71476
rect 256068 71466 256096 73630
rect 269396 72072 269448 72078
rect 269396 72014 269448 72020
rect 269408 71602 269436 72014
rect 270328 71602 270356 82418
rect 269396 71596 269448 71602
rect 269396 71538 269448 71544
rect 270316 71596 270368 71602
rect 270316 71538 270368 71544
rect 256056 71460 256108 71466
rect 256056 71402 256108 71408
rect 111800 71392 111852 71398
rect 111800 71334 111852 71340
rect 270604 3670 270632 350775
rect 270696 333713 270724 700062
rect 270776 699984 270828 699990
rect 270776 699926 270828 699932
rect 270682 333704 270738 333713
rect 270682 333639 270738 333648
rect 270788 317801 270816 699926
rect 270880 342689 270908 700198
rect 271144 586560 271196 586566
rect 271144 586502 271196 586508
rect 271156 586090 271184 586502
rect 272248 586492 272300 586498
rect 272248 586434 272300 586440
rect 271144 586084 271196 586090
rect 271144 586026 271196 586032
rect 272156 511556 272208 511562
rect 272156 511498 272208 511504
rect 271052 382696 271104 382702
rect 271052 382638 271104 382644
rect 270960 382492 271012 382498
rect 270960 382434 271012 382440
rect 270972 382158 271000 382434
rect 270960 382152 271012 382158
rect 270960 382094 271012 382100
rect 271064 382022 271092 382638
rect 271972 382492 272024 382498
rect 271972 382434 272024 382440
rect 271052 382016 271104 382022
rect 271052 381958 271104 381964
rect 271512 357876 271564 357882
rect 271512 357818 271564 357824
rect 270866 342680 270922 342689
rect 270866 342615 270922 342624
rect 270774 317792 270830 317801
rect 270774 317727 270830 317736
rect 271524 71738 271552 357818
rect 271984 313274 272012 382434
rect 272064 382016 272116 382022
rect 272064 381958 272116 381964
rect 271972 313268 272024 313274
rect 271972 313210 272024 313216
rect 272076 313206 272104 381958
rect 272168 316266 272196 511498
rect 272156 316260 272208 316266
rect 272156 316202 272208 316208
rect 272260 313410 272288 586434
rect 272614 327584 272670 327593
rect 272996 327570 273024 700266
rect 364996 700262 365024 703520
rect 397472 700670 397500 703520
rect 397460 700664 397512 700670
rect 397460 700606 397512 700612
rect 364984 700256 365036 700262
rect 364984 700198 365036 700204
rect 312084 700188 312136 700194
rect 312084 700130 312136 700136
rect 306196 586560 306248 586566
rect 306196 586502 306248 586508
rect 292948 586424 293000 586430
rect 292948 586366 293000 586372
rect 300216 586424 300268 586430
rect 300216 586366 300268 586372
rect 292960 586158 292988 586366
rect 292948 586152 293000 586158
rect 292948 586094 293000 586100
rect 294328 586152 294380 586158
rect 294328 586094 294380 586100
rect 288532 585948 288584 585954
rect 288532 585890 288584 585896
rect 275928 582344 275980 582350
rect 275928 582286 275980 582292
rect 275940 580718 275968 582286
rect 275928 580712 275980 580718
rect 275928 580654 275980 580660
rect 273812 569628 273864 569634
rect 273812 569570 273864 569576
rect 273824 565894 273852 569570
rect 273812 565888 273864 565894
rect 273812 565830 273864 565836
rect 275284 565888 275336 565894
rect 275284 565830 275336 565836
rect 275296 562834 275324 565830
rect 275284 562828 275336 562834
rect 275284 562770 275336 562776
rect 275284 382696 275336 382702
rect 275284 382638 275336 382644
rect 275296 382362 275324 382638
rect 275192 382356 275244 382362
rect 275192 382298 275244 382304
rect 275284 382356 275336 382362
rect 275284 382298 275336 382304
rect 275204 381954 275232 382298
rect 275192 381948 275244 381954
rect 275192 381890 275244 381896
rect 273168 359440 273220 359446
rect 273168 359382 273220 359388
rect 272670 327542 273024 327570
rect 272614 327519 272670 327528
rect 272248 313404 272300 313410
rect 272248 313346 272300 313352
rect 272064 313200 272116 313206
rect 272064 313142 272116 313148
rect 273180 276010 273208 359382
rect 273352 359372 273404 359378
rect 273352 359314 273404 359320
rect 273260 356312 273312 356318
rect 273260 356254 273312 356260
rect 273168 276004 273220 276010
rect 273168 275946 273220 275952
rect 273272 272134 273300 356254
rect 273260 272128 273312 272134
rect 273260 272070 273312 272076
rect 273364 130626 273392 359314
rect 273444 359236 273496 359242
rect 273444 359178 273496 359184
rect 273352 130620 273404 130626
rect 273352 130562 273404 130568
rect 273364 130286 273392 130562
rect 273352 130280 273404 130286
rect 273352 130222 273404 130228
rect 273456 72010 273484 359178
rect 274364 358420 274416 358426
rect 274364 358362 274416 358368
rect 274376 355436 274404 358362
rect 275940 356318 275968 580654
rect 279608 562828 279660 562834
rect 279608 562770 279660 562776
rect 279620 559314 279648 562770
rect 279620 559286 279740 559314
rect 279712 556510 279740 559286
rect 279700 556504 279752 556510
rect 279700 556446 279752 556452
rect 285496 556436 285548 556442
rect 285496 556378 285548 556384
rect 285508 549778 285536 556378
rect 285496 549772 285548 549778
rect 285496 549714 285548 549720
rect 286232 440156 286284 440162
rect 286232 440098 286284 440104
rect 286244 386306 286272 440098
rect 278136 386300 278188 386306
rect 278136 386242 278188 386248
rect 286232 386300 286284 386306
rect 286232 386242 286284 386248
rect 278148 386209 278176 386242
rect 278134 386200 278190 386209
rect 278134 386135 278190 386144
rect 278228 382424 278280 382430
rect 278228 382366 278280 382372
rect 279516 382424 279568 382430
rect 279516 382366 279568 382372
rect 279700 382424 279752 382430
rect 279700 382366 279752 382372
rect 278240 373810 278268 382366
rect 279528 382158 279556 382366
rect 279712 382294 279740 382366
rect 279700 382288 279752 382294
rect 279700 382230 279752 382236
rect 279516 382152 279568 382158
rect 279516 382094 279568 382100
rect 278240 373782 278360 373810
rect 278332 363610 278360 373782
rect 278332 363582 278544 363610
rect 278516 359242 278544 363582
rect 278596 359440 278648 359446
rect 278596 359382 278648 359388
rect 278608 359242 278636 359382
rect 278504 359236 278556 359242
rect 278504 359178 278556 359184
rect 278596 359236 278648 359242
rect 278596 359178 278648 359184
rect 275928 356312 275980 356318
rect 275928 356254 275980 356260
rect 275940 355586 275968 356254
rect 275940 355558 276244 355586
rect 276216 355450 276244 355558
rect 278516 355450 278544 359178
rect 276216 355422 276598 355450
rect 278516 355422 278622 355450
rect 279712 354890 279740 382230
rect 286244 359378 286272 386242
rect 286324 382696 286376 382702
rect 286324 382638 286376 382644
rect 286336 382294 286364 382638
rect 286324 382288 286376 382294
rect 286324 382230 286376 382236
rect 288544 373810 288572 585890
rect 290648 549772 290700 549778
rect 290648 549714 290700 549720
rect 290660 540258 290688 549714
rect 290648 540252 290700 540258
rect 290648 540194 290700 540200
rect 293316 540184 293368 540190
rect 293316 540126 293368 540132
rect 293328 537266 293356 540126
rect 293316 537260 293368 537266
rect 293316 537202 293368 537208
rect 291384 386368 291436 386374
rect 291384 386310 291436 386316
rect 291396 386170 291424 386310
rect 291384 386164 291436 386170
rect 291384 386106 291436 386112
rect 288544 373782 288664 373810
rect 288636 363610 288664 373782
rect 288636 363582 288848 363610
rect 286232 359372 286284 359378
rect 286232 359314 286284 359320
rect 282644 358420 282696 358426
rect 282644 358362 282696 358368
rect 282656 355436 282684 358362
rect 284668 357808 284720 357814
rect 284668 357750 284720 357756
rect 284680 355436 284708 357750
rect 286244 355450 286272 359314
rect 288820 359242 288848 363582
rect 294340 359242 294368 586094
rect 294420 537260 294472 537266
rect 294420 537202 294472 537208
rect 294432 534410 294460 537202
rect 294420 534404 294472 534410
rect 294420 534346 294472 534352
rect 298008 534268 298060 534274
rect 298008 534210 298060 534216
rect 298020 524006 298048 534210
rect 298836 529916 298888 529922
rect 298836 529858 298888 529864
rect 298848 527082 298876 529858
rect 298756 527054 298876 527082
rect 298008 524000 298060 524006
rect 298008 523942 298060 523948
rect 298756 522646 298784 527054
rect 300124 524000 300176 524006
rect 300124 523942 300176 523948
rect 295064 522640 295116 522646
rect 295064 522582 295116 522588
rect 298744 522640 298796 522646
rect 298744 522582 298796 522588
rect 295076 511562 295104 522582
rect 300136 519110 300164 523942
rect 300124 519104 300176 519110
rect 300124 519046 300176 519052
rect 295064 511556 295116 511562
rect 295064 511498 295116 511504
rect 298834 386472 298890 386481
rect 298744 386436 298796 386442
rect 298834 386407 298836 386416
rect 298744 386378 298796 386384
rect 298888 386407 298890 386416
rect 298836 386378 298888 386384
rect 298756 386170 298784 386378
rect 298744 386164 298796 386170
rect 298744 386106 298796 386112
rect 295892 382288 295944 382294
rect 295892 382230 295944 382236
rect 295904 381954 295932 382230
rect 295892 381948 295944 381954
rect 295892 381890 295944 381896
rect 288808 359236 288860 359242
rect 288808 359178 288860 359184
rect 292948 359236 293000 359242
rect 292948 359178 293000 359184
rect 294328 359236 294380 359242
rect 294328 359178 294380 359184
rect 288820 355450 288848 359178
rect 290924 357808 290976 357814
rect 290924 357750 290976 357756
rect 286244 355422 286718 355450
rect 288820 355422 288926 355450
rect 290936 355436 290964 357750
rect 292960 355436 292988 359178
rect 294972 358488 295024 358494
rect 294972 358430 295024 358436
rect 294984 355436 295012 358430
rect 300228 358358 300256 586366
rect 306208 586226 306236 586502
rect 306196 586220 306248 586226
rect 306196 586162 306248 586168
rect 309784 559360 309836 559366
rect 309784 559302 309836 559308
rect 309796 544610 309824 559302
rect 307668 544604 307720 544610
rect 307668 544546 307720 544552
rect 309784 544604 309836 544610
rect 309784 544546 309836 544552
rect 307680 536586 307708 544546
rect 304724 536580 304776 536586
rect 304724 536522 304776 536528
rect 307668 536580 307720 536586
rect 307668 536522 307720 536528
rect 304736 534546 304764 536522
rect 303252 534540 303304 534546
rect 303252 534482 303304 534488
rect 304724 534540 304776 534546
rect 304724 534482 304776 534488
rect 303264 529990 303292 534482
rect 303252 529984 303304 529990
rect 303252 529926 303304 529932
rect 301596 519104 301648 519110
rect 301596 519046 301648 519052
rect 301608 516730 301636 519046
rect 301596 516724 301648 516730
rect 301596 516666 301648 516672
rect 303160 516724 303212 516730
rect 303160 516666 303212 516672
rect 303172 515234 303200 516666
rect 303160 515228 303212 515234
rect 303160 515170 303212 515176
rect 307392 515160 307444 515166
rect 307392 515102 307444 515108
rect 307404 509726 307432 515102
rect 307392 509720 307444 509726
rect 307392 509662 307444 509668
rect 307404 487286 307432 509662
rect 307392 487280 307444 487286
rect 307392 487222 307444 487228
rect 307576 487280 307628 487286
rect 307576 487222 307628 487228
rect 307588 476898 307616 487222
rect 307404 476870 307616 476898
rect 307404 466682 307432 476870
rect 307392 466676 307444 466682
rect 307392 466618 307444 466624
rect 307576 466676 307628 466682
rect 307576 466618 307628 466624
rect 307588 466562 307616 466618
rect 307404 466534 307616 466562
rect 307404 446078 307432 466534
rect 307392 446072 307444 446078
rect 307392 446014 307444 446020
rect 307576 446072 307628 446078
rect 307576 446014 307628 446020
rect 307588 435690 307616 446014
rect 307404 435662 307616 435690
rect 307404 425474 307432 435662
rect 307392 425468 307444 425474
rect 307392 425410 307444 425416
rect 307576 425468 307628 425474
rect 307576 425410 307628 425416
rect 307588 425354 307616 425410
rect 307404 425326 307616 425354
rect 303896 404864 303948 404870
rect 303896 404806 303948 404812
rect 307404 404818 307432 425326
rect 303908 384946 303936 404806
rect 307404 404790 307616 404818
rect 307588 394482 307616 404790
rect 307404 394454 307616 394482
rect 303896 384940 303948 384946
rect 303896 384882 303948 384888
rect 307404 384266 307432 394454
rect 309046 386472 309102 386481
rect 309046 386407 309102 386416
rect 309060 386374 309088 386407
rect 309048 386368 309100 386374
rect 309048 386310 309100 386316
rect 307392 384260 307444 384266
rect 307392 384202 307444 384208
rect 307576 384260 307628 384266
rect 307576 384202 307628 384208
rect 307588 384146 307616 384202
rect 307404 384118 307616 384146
rect 301688 382696 301740 382702
rect 301688 382638 301740 382644
rect 301700 382090 301728 382638
rect 301688 382084 301740 382090
rect 301688 382026 301740 382032
rect 301700 359378 301728 382026
rect 307404 363610 307432 384118
rect 307404 363582 307616 363610
rect 306932 359440 306984 359446
rect 306932 359382 306984 359388
rect 307024 359440 307076 359446
rect 307024 359382 307076 359388
rect 301228 359372 301280 359378
rect 301228 359314 301280 359320
rect 301688 359372 301740 359378
rect 301688 359314 301740 359320
rect 299020 358352 299072 358358
rect 299020 358294 299072 358300
rect 300216 358352 300268 358358
rect 300216 358294 300268 358300
rect 296996 357876 297048 357882
rect 296996 357818 297048 357824
rect 297008 355436 297036 357818
rect 299032 355436 299060 358294
rect 301240 355436 301268 359314
rect 306944 359310 306972 359382
rect 306932 359304 306984 359310
rect 306932 359246 306984 359252
rect 307036 359242 307064 359382
rect 307588 359242 307616 363582
rect 307024 359236 307076 359242
rect 307024 359178 307076 359184
rect 307576 359236 307628 359242
rect 307576 359178 307628 359184
rect 305276 358556 305328 358562
rect 305276 358498 305328 358504
rect 303252 358488 303304 358494
rect 303252 358430 303304 358436
rect 303264 355436 303292 358430
rect 305288 355436 305316 358498
rect 307588 355450 307616 359178
rect 311348 357944 311400 357950
rect 311348 357886 311400 357892
rect 309324 357740 309376 357746
rect 309324 357682 309376 357688
rect 307326 355422 307616 355450
rect 309336 355436 309364 357682
rect 311360 355436 311388 357886
rect 280264 354890 280646 354906
rect 273536 354884 273588 354890
rect 273536 354826 273588 354832
rect 279700 354884 279752 354890
rect 279700 354826 279752 354832
rect 280252 354884 280646 354890
rect 280304 354878 280646 354884
rect 280252 354826 280304 354832
rect 272340 72004 272392 72010
rect 272340 71946 272392 71952
rect 273444 72004 273496 72010
rect 273444 71946 273496 71952
rect 271512 71732 271564 71738
rect 271512 71674 271564 71680
rect 272352 71670 272380 71946
rect 273548 71738 273576 354826
rect 311532 354136 311584 354142
rect 311532 354078 311584 354084
rect 311544 352073 311572 354078
rect 311530 352064 311586 352073
rect 311530 351999 311586 352008
rect 312096 318753 312124 700130
rect 429856 700126 429884 703520
rect 462332 700670 462360 703520
rect 462320 700664 462372 700670
rect 462320 700606 462372 700612
rect 429844 700120 429896 700126
rect 429844 700062 429896 700068
rect 494808 700058 494836 703520
rect 527192 700670 527220 703520
rect 527180 700664 527232 700670
rect 527180 700606 527232 700612
rect 312176 700052 312228 700058
rect 312176 699994 312228 700000
rect 312728 700052 312780 700058
rect 312728 699994 312780 700000
rect 494796 700052 494848 700058
rect 494796 699994 494848 700000
rect 312188 325009 312216 699994
rect 312360 586288 312412 586294
rect 312360 586230 312412 586236
rect 312268 359304 312320 359310
rect 312268 359246 312320 359252
rect 312174 325000 312230 325009
rect 312174 324935 312230 324944
rect 312082 318744 312138 318753
rect 312082 318679 312138 318688
rect 310638 316266 310928 316282
rect 275284 316260 275336 316266
rect 310638 316260 310940 316266
rect 310638 316254 310888 316260
rect 275284 316202 275336 316208
rect 310888 316202 310940 316208
rect 275296 315602 275324 316202
rect 294262 315846 294460 315874
rect 273640 313342 273668 315588
rect 275296 315574 275968 315602
rect 273628 313336 273680 313342
rect 273628 313278 273680 313284
rect 275940 272270 275968 315574
rect 277688 313342 277716 315588
rect 279712 315574 279910 315602
rect 277676 313336 277728 313342
rect 277676 313278 277728 313284
rect 279712 313206 279740 315574
rect 281920 313274 281948 315588
rect 283944 313410 283972 315588
rect 285968 313478 285996 315588
rect 287992 313478 288020 315588
rect 285956 313472 286008 313478
rect 285956 313414 286008 313420
rect 287980 313472 288032 313478
rect 287980 313414 288032 313420
rect 283932 313404 283984 313410
rect 283932 313346 283984 313352
rect 281908 313268 281960 313274
rect 281908 313210 281960 313216
rect 279700 313200 279752 313206
rect 279700 313142 279752 313148
rect 275928 272264 275980 272270
rect 275928 272206 275980 272212
rect 275940 202842 275968 272206
rect 276664 272128 276716 272134
rect 276664 272070 276716 272076
rect 276676 270842 276704 272070
rect 276664 270836 276716 270842
rect 276664 270778 276716 270784
rect 275928 202836 275980 202842
rect 275928 202778 275980 202784
rect 279712 72078 279740 313142
rect 281920 312118 281948 313210
rect 283944 312118 283972 313346
rect 290016 312934 290044 315588
rect 292224 313410 292252 315588
rect 292212 313404 292264 313410
rect 292212 313346 292264 313352
rect 290004 312928 290056 312934
rect 290004 312870 290056 312876
rect 294432 312338 294460 315846
rect 296272 313274 296300 315588
rect 298310 315574 298784 315602
rect 296260 313268 296312 313274
rect 296260 313210 296312 313216
rect 297272 313268 297324 313274
rect 297272 313210 297324 313216
rect 294340 312310 294460 312338
rect 281172 312112 281224 312118
rect 281172 312054 281224 312060
rect 281908 312112 281960 312118
rect 281908 312054 281960 312060
rect 282644 312112 282696 312118
rect 282644 312054 282696 312060
rect 283932 312112 283984 312118
rect 283932 312054 283984 312060
rect 279700 72072 279752 72078
rect 279700 72014 279752 72020
rect 280160 72072 280212 72078
rect 280160 72014 280212 72020
rect 272432 71732 272484 71738
rect 272432 71674 272484 71680
rect 273536 71732 273588 71738
rect 273536 71674 273588 71680
rect 272340 71664 272392 71670
rect 272340 71606 272392 71612
rect 272444 71398 272472 71674
rect 280172 71466 280200 72014
rect 281184 71942 281212 312054
rect 282656 276486 282684 312054
rect 285588 276616 285640 276622
rect 285588 276558 285640 276564
rect 282644 276480 282696 276486
rect 282644 276422 282696 276428
rect 282656 276282 282684 276422
rect 285600 276350 285628 276558
rect 294340 276418 294368 312310
rect 295800 276616 295852 276622
rect 295800 276558 295852 276564
rect 294328 276412 294380 276418
rect 294328 276354 294380 276360
rect 285588 276344 285640 276350
rect 285588 276286 285640 276292
rect 295812 276282 295840 276558
rect 282644 276276 282696 276282
rect 282644 276218 282696 276224
rect 295800 276276 295852 276282
rect 295800 276218 295852 276224
rect 291476 130280 291528 130286
rect 291476 130222 291528 130228
rect 291488 125594 291516 130222
rect 291476 125588 291528 125594
rect 291476 125530 291528 125536
rect 293592 125588 293644 125594
rect 293592 125530 293644 125536
rect 293604 116278 293632 125530
rect 293592 116272 293644 116278
rect 293592 116214 293644 116220
rect 294696 116272 294748 116278
rect 294696 116214 294748 116220
rect 294708 114782 294736 116214
rect 294696 114776 294748 114782
rect 294696 114718 294748 114724
rect 296444 114776 296496 114782
rect 296444 114718 296496 114724
rect 296456 111858 296484 114718
rect 296444 111852 296496 111858
rect 296444 111794 296496 111800
rect 297284 71942 297312 313210
rect 298756 313206 298784 315574
rect 298744 313200 298796 313206
rect 298744 313142 298796 313148
rect 298756 276282 298784 313142
rect 300320 312866 300348 315588
rect 300308 312860 300360 312866
rect 300308 312802 300360 312808
rect 302528 312798 302556 315588
rect 302516 312792 302568 312798
rect 302516 312734 302568 312740
rect 304552 312050 304580 315588
rect 306576 313070 306604 315588
rect 308600 313546 308628 315588
rect 308588 313540 308640 313546
rect 308588 313482 308640 313488
rect 306564 313064 306616 313070
rect 306564 313006 306616 313012
rect 307576 313064 307628 313070
rect 307576 313006 307628 313012
rect 303896 312044 303948 312050
rect 303896 311986 303948 311992
rect 304540 312044 304592 312050
rect 304540 311986 304592 311992
rect 298744 276276 298796 276282
rect 298744 276218 298796 276224
rect 297364 111852 297416 111858
rect 297364 111794 297416 111800
rect 297376 109342 297404 111794
rect 297364 109336 297416 109342
rect 297364 109278 297416 109284
rect 300216 109336 300268 109342
rect 300216 109278 300268 109284
rect 300228 107386 300256 109278
rect 300228 107358 300348 107386
rect 300320 101590 300348 107358
rect 300308 101584 300360 101590
rect 300308 101526 300360 101532
rect 301780 101584 301832 101590
rect 301780 101526 301832 101532
rect 301792 94246 301820 101526
rect 303908 94926 303936 311986
rect 307588 276622 307616 313006
rect 307024 276616 307076 276622
rect 307024 276558 307076 276564
rect 307576 276616 307628 276622
rect 307576 276558 307628 276564
rect 306196 276276 306248 276282
rect 306196 276218 306248 276224
rect 306208 275942 306236 276218
rect 307036 276078 307064 276558
rect 312084 276548 312136 276554
rect 312084 276490 312136 276496
rect 312096 276078 312124 276490
rect 307024 276072 307076 276078
rect 307024 276014 307076 276020
rect 312084 276072 312136 276078
rect 312084 276014 312136 276020
rect 306196 275936 306248 275942
rect 306196 275878 306248 275884
rect 303896 94920 303948 94926
rect 303896 94862 303948 94868
rect 301780 94240 301832 94246
rect 301780 94182 301832 94188
rect 303908 75954 303936 94862
rect 304724 94172 304776 94178
rect 304724 94114 304776 94120
rect 304736 90438 304764 94114
rect 304724 90432 304776 90438
rect 304724 90374 304776 90380
rect 307668 90432 307720 90438
rect 307668 90374 307720 90380
rect 307680 86902 307708 90374
rect 307668 86896 307720 86902
rect 307668 86838 307720 86844
rect 312084 86828 312136 86834
rect 312084 86770 312136 86776
rect 312096 81190 312124 86770
rect 312084 81184 312136 81190
rect 312084 81126 312136 81132
rect 303896 75948 303948 75954
rect 303896 75890 303948 75896
rect 312280 74338 312308 359246
rect 312372 342961 312400 586230
rect 312636 384940 312688 384946
rect 312636 384882 312688 384888
rect 312544 359440 312596 359446
rect 312544 359382 312596 359388
rect 312452 359236 312504 359242
rect 312452 359178 312504 359184
rect 312358 342952 312414 342961
rect 312358 342887 312414 342896
rect 312464 275210 312492 359178
rect 312556 276554 312584 359382
rect 312648 312050 312676 384882
rect 312740 316266 312768 699994
rect 527192 699922 527220 700606
rect 559668 699990 559696 703520
rect 559656 699984 559708 699990
rect 559656 699926 559708 699932
rect 314476 699916 314528 699922
rect 314476 699858 314528 699864
rect 527180 699916 527232 699922
rect 527180 699858 527232 699864
rect 579896 699916 579948 699922
rect 579896 699858 579948 699864
rect 313740 586628 313792 586634
rect 313740 586570 313792 586576
rect 313752 586362 313780 586570
rect 313648 586356 313700 586362
rect 313648 586298 313700 586304
rect 313740 586356 313792 586362
rect 313740 586298 313792 586304
rect 312820 586288 312872 586294
rect 312820 586230 312872 586236
rect 312728 316260 312780 316266
rect 312728 316202 312780 316208
rect 312832 313342 312860 586230
rect 313660 586022 313688 586298
rect 313648 586016 313700 586022
rect 313648 585958 313700 585964
rect 313556 382628 313608 382634
rect 313556 382570 313608 382576
rect 313568 382090 313596 382570
rect 313556 382084 313608 382090
rect 313556 382026 313608 382032
rect 313556 354000 313608 354006
rect 313556 353942 313608 353948
rect 313568 339969 313596 353942
rect 313554 339960 313610 339969
rect 313554 339895 313610 339904
rect 313554 328264 313610 328273
rect 313554 328199 313610 328208
rect 313568 327593 313596 328199
rect 313554 327584 313610 327593
rect 313554 327519 313610 327528
rect 312820 313336 312872 313342
rect 312820 313278 312872 313284
rect 312636 312044 312688 312050
rect 312636 311986 312688 311992
rect 312544 276548 312596 276554
rect 312544 276490 312596 276496
rect 312464 275182 312584 275210
rect 312556 272066 312584 275182
rect 312544 272060 312596 272066
rect 312544 272002 312596 272008
rect 312556 265010 312584 272002
rect 312556 264982 312768 265010
rect 312740 200190 312768 264982
rect 312728 200184 312780 200190
rect 312728 200126 312780 200132
rect 312280 74310 312400 74338
rect 312372 72146 312400 74310
rect 313568 72146 313596 327519
rect 313660 313206 313688 585958
rect 313648 313200 313700 313206
rect 313648 313142 313700 313148
rect 313752 313070 313780 586298
rect 314292 582276 314344 582282
rect 314292 582218 314344 582224
rect 314200 547596 314252 547602
rect 314200 547538 314252 547544
rect 314016 385756 314068 385762
rect 314016 385698 314068 385704
rect 313924 382084 313976 382090
rect 313924 382026 313976 382032
rect 313832 381948 313884 381954
rect 313832 381890 313884 381896
rect 313844 328273 313872 381890
rect 313830 328264 313886 328273
rect 313830 328199 313886 328208
rect 313936 313274 313964 382026
rect 314028 345817 314056 385698
rect 314108 382220 314160 382226
rect 314108 382162 314160 382168
rect 314014 345808 314070 345817
rect 314014 345743 314070 345752
rect 314028 344593 314056 345743
rect 314014 344584 314070 344593
rect 314014 344519 314070 344528
rect 314016 334144 314068 334150
rect 314016 334086 314068 334092
rect 314028 333849 314056 334086
rect 314014 333840 314070 333849
rect 314014 333775 314070 333784
rect 314016 333464 314068 333470
rect 314016 333406 314068 333412
rect 313924 313268 313976 313274
rect 313924 313210 313976 313216
rect 313740 313064 313792 313070
rect 313740 313006 313792 313012
rect 314028 271998 314056 333406
rect 314120 330993 314148 382162
rect 314212 348809 314240 547538
rect 314304 544950 314332 582218
rect 314292 544944 314344 544950
rect 314292 544886 314344 544892
rect 314198 348800 314254 348809
rect 314198 348735 314254 348744
rect 314198 344584 314254 344593
rect 314198 344519 314254 344528
rect 314106 330984 314162 330993
rect 314106 330919 314162 330928
rect 314016 271992 314068 271998
rect 314016 271934 314068 271940
rect 314028 270910 314056 271934
rect 314016 270904 314068 270910
rect 314016 270846 314068 270852
rect 312360 72140 312412 72146
rect 312360 72082 312412 72088
rect 313556 72140 313608 72146
rect 313556 72082 313608 72088
rect 281172 71936 281224 71942
rect 281172 71878 281224 71884
rect 297272 71936 297324 71942
rect 297272 71878 297324 71884
rect 281184 71670 281212 71878
rect 281172 71664 281224 71670
rect 281172 71606 281224 71612
rect 297284 71534 297312 71878
rect 312372 71534 312400 72082
rect 313568 71806 313596 72082
rect 314120 71874 314148 330919
rect 314212 92410 314240 344519
rect 314304 336569 314332 544886
rect 314382 402248 314438 402257
rect 314382 402183 314438 402192
rect 314396 386374 314424 402183
rect 314384 386368 314436 386374
rect 314384 386310 314436 386316
rect 314396 385762 314424 386310
rect 314384 385756 314436 385762
rect 314384 385698 314436 385704
rect 314382 348800 314438 348809
rect 314382 348735 314438 348744
rect 314290 336560 314346 336569
rect 314290 336495 314346 336504
rect 314304 333470 314332 336495
rect 314292 333464 314344 333470
rect 314292 333406 314344 333412
rect 314396 272406 314424 348735
rect 314488 322017 314516 699858
rect 579908 698057 579936 699858
rect 579894 698048 579950 698057
rect 579894 697983 579950 697992
rect 578514 674656 578570 674665
rect 578514 674591 578570 674600
rect 578528 674218 578556 674591
rect 561496 674212 561548 674218
rect 561496 674154 561548 674160
rect 578516 674212 578568 674218
rect 578516 674154 578568 674160
rect 316408 586560 316460 586566
rect 316408 586502 316460 586508
rect 326896 586560 326948 586566
rect 326896 586502 326948 586508
rect 337016 586560 337068 586566
rect 337016 586502 337068 586508
rect 347412 586560 347464 586566
rect 347412 586502 347464 586508
rect 357624 586560 357676 586566
rect 357624 586502 357676 586508
rect 463698 586528 463754 586537
rect 316420 586226 316448 586502
rect 326908 586226 326936 586502
rect 337028 586226 337056 586502
rect 341524 586356 341576 586362
rect 341524 586298 341576 586304
rect 316408 586220 316460 586226
rect 316408 586162 316460 586168
rect 326896 586220 326948 586226
rect 326896 586162 326948 586168
rect 337016 586220 337068 586226
rect 337016 586162 337068 586168
rect 341536 583930 341564 586298
rect 347424 586226 347452 586502
rect 357636 586226 357664 586502
rect 365444 586492 365496 586498
rect 365444 586434 365496 586440
rect 368020 586492 368072 586498
rect 368020 586434 368072 586440
rect 378232 586492 378284 586498
rect 378232 586434 378284 586440
rect 388628 586492 388680 586498
rect 388628 586434 388680 586440
rect 398840 586492 398892 586498
rect 398840 586434 398892 586440
rect 409236 586492 409288 586498
rect 409236 586434 409288 586440
rect 415124 586492 415176 586498
rect 463698 586463 463700 586472
rect 415124 586434 415176 586440
rect 463752 586463 463754 586472
rect 473910 586528 473966 586537
rect 473910 586463 473966 586472
rect 485780 586492 485832 586498
rect 463700 586434 463752 586440
rect 347412 586220 347464 586226
rect 347412 586162 347464 586168
rect 357624 586220 357676 586226
rect 357624 586162 357676 586168
rect 365456 583930 365484 586434
rect 368032 586226 368060 586434
rect 378244 586226 378272 586434
rect 388640 586226 388668 586434
rect 398852 586226 398880 586434
rect 409248 586226 409276 586434
rect 415136 586294 415164 586434
rect 473924 586430 473952 586463
rect 485780 586434 485832 586440
rect 437756 586424 437808 586430
rect 456248 586424 456300 586430
rect 437756 586366 437808 586372
rect 413652 586288 413704 586294
rect 413652 586230 413704 586236
rect 415124 586288 415176 586294
rect 415124 586230 415176 586236
rect 432786 586256 432842 586265
rect 368020 586220 368072 586226
rect 368020 586162 368072 586168
rect 378232 586220 378284 586226
rect 378232 586162 378284 586168
rect 388628 586220 388680 586226
rect 388628 586162 388680 586168
rect 398840 586220 398892 586226
rect 398840 586162 398892 586168
rect 409236 586220 409288 586226
rect 409236 586162 409288 586168
rect 413664 583930 413692 586230
rect 432786 586191 432788 586200
rect 432840 586191 432842 586200
rect 432788 586162 432840 586168
rect 437768 583930 437796 586366
rect 442920 586350 443040 586378
rect 456340 586424 456392 586430
rect 456300 586372 456340 586378
rect 456248 586366 456392 586372
rect 473912 586424 473964 586430
rect 473912 586366 473964 586372
rect 476856 586424 476908 586430
rect 476948 586424 477000 586430
rect 476908 586372 476948 586378
rect 476856 586366 477000 586372
rect 456260 586350 456380 586366
rect 476868 586350 476988 586366
rect 442920 586265 442948 586350
rect 443012 586294 443040 586350
rect 443000 586288 443052 586294
rect 442906 586256 442962 586265
rect 443000 586230 443052 586236
rect 442906 586191 442962 586200
rect 461676 586016 461728 586022
rect 461676 585958 461728 585964
rect 461688 583930 461716 585958
rect 485792 583930 485820 586434
rect 533988 586152 534040 586158
rect 533988 586094 534040 586100
rect 509884 586084 509936 586090
rect 509884 586026 509936 586032
rect 509896 583930 509924 586026
rect 534000 583930 534028 586094
rect 557908 585948 557960 585954
rect 557908 585890 557960 585896
rect 557920 583930 557948 585890
rect 341536 583902 341826 583930
rect 365456 583902 365746 583930
rect 413664 583902 413954 583930
rect 437768 583902 438058 583930
rect 461688 583902 461978 583930
rect 485792 583902 486082 583930
rect 509896 583902 510186 583930
rect 534000 583902 534290 583930
rect 557920 583902 558210 583930
rect 318616 582956 318668 582962
rect 318616 582898 318668 582904
rect 560852 582956 560904 582962
rect 560852 582898 560904 582904
rect 315028 580712 315080 580718
rect 315026 580680 315028 580689
rect 315080 580680 315082 580689
rect 315026 580615 315082 580624
rect 317972 576292 318024 576298
rect 317972 576234 318024 576240
rect 317984 572694 318012 576234
rect 317144 572688 317196 572694
rect 317144 572630 317196 572636
rect 317972 572688 318024 572694
rect 317972 572630 318024 572636
rect 317156 562358 317184 572630
rect 315028 562352 315080 562358
rect 315028 562294 315080 562300
rect 317144 562352 317196 562358
rect 317144 562294 317196 562300
rect 315040 559434 315068 562294
rect 315028 559428 315080 559434
rect 315028 559370 315080 559376
rect 318628 547602 318656 582898
rect 319444 582276 319496 582282
rect 319444 582218 319496 582224
rect 558460 582276 558512 582282
rect 558460 582218 558512 582224
rect 319456 576298 319484 582218
rect 319444 576292 319496 576298
rect 319444 576234 319496 576240
rect 318616 547596 318668 547602
rect 318616 547538 318668 547544
rect 315028 544944 315080 544950
rect 315026 544912 315028 544921
rect 315080 544912 315082 544921
rect 315026 544847 315082 544856
rect 558472 512174 558500 582218
rect 560864 547777 560892 582898
rect 560850 547768 560906 547777
rect 560850 547703 560906 547712
rect 558460 512168 558512 512174
rect 558460 512110 558512 512116
rect 558920 512168 558972 512174
rect 558920 512110 558972 512116
rect 558932 512077 558960 512110
rect 558918 512068 558974 512077
rect 558918 512003 558974 512012
rect 315028 509720 315080 509726
rect 315026 509688 315028 509697
rect 315080 509688 315082 509697
rect 315026 509623 315082 509632
rect 315026 473104 315082 473113
rect 315026 473039 315082 473048
rect 315040 472598 315068 473039
rect 315028 472592 315080 472598
rect 315028 472534 315080 472540
rect 558918 440804 558974 440813
rect 558918 440739 558974 440748
rect 558932 440502 558960 440739
rect 558460 440496 558512 440502
rect 558460 440438 558512 440444
rect 558920 440496 558972 440502
rect 558920 440438 558972 440444
rect 558472 386306 558500 440438
rect 560850 405376 560906 405385
rect 560850 405311 560906 405320
rect 558460 386300 558512 386306
rect 558460 386242 558512 386248
rect 560864 384946 560892 405311
rect 560852 384940 560904 384946
rect 560852 384882 560904 384888
rect 331508 382702 331536 383996
rect 331496 382696 331548 382702
rect 331496 382638 331548 382644
rect 355612 382566 355640 383996
rect 355600 382560 355652 382566
rect 355600 382502 355652 382508
rect 379532 382498 379560 383996
rect 379520 382492 379572 382498
rect 379520 382434 379572 382440
rect 403636 382430 403664 383996
rect 403624 382424 403676 382430
rect 403624 382366 403676 382372
rect 316408 382288 316460 382294
rect 316408 382230 316460 382236
rect 316420 381954 316448 382230
rect 427740 382226 427768 383996
rect 475948 382294 475976 383996
rect 475936 382288 475988 382294
rect 475936 382230 475988 382236
rect 427728 382220 427780 382226
rect 427728 382162 427780 382168
rect 499868 382158 499896 383996
rect 499856 382152 499908 382158
rect 499856 382094 499908 382100
rect 523972 382090 524000 383996
rect 523960 382084 524012 382090
rect 523960 382026 524012 382032
rect 548076 382022 548104 383996
rect 548064 382016 548116 382022
rect 548064 381958 548116 381964
rect 316408 381948 316460 381954
rect 316408 381890 316460 381896
rect 317144 357808 317196 357814
rect 317144 357750 317196 357756
rect 315672 357740 315724 357746
rect 315672 357682 315724 357688
rect 314474 322008 314530 322017
rect 314474 321943 314530 321952
rect 314384 272400 314436 272406
rect 314384 272342 314436 272348
rect 314292 270904 314344 270910
rect 314292 270846 314344 270852
rect 314304 234705 314332 270846
rect 314396 238474 314424 272342
rect 315028 270836 315080 270842
rect 315028 270778 315080 270784
rect 315040 270337 315068 270778
rect 315026 270328 315082 270337
rect 315026 270263 315082 270272
rect 314384 238468 314436 238474
rect 314384 238410 314436 238416
rect 314290 234696 314346 234705
rect 314290 234631 314346 234640
rect 315028 200184 315080 200190
rect 315028 200126 315080 200132
rect 315040 199073 315068 200126
rect 315026 199064 315082 199073
rect 315026 198999 315082 199008
rect 315684 163441 315712 357682
rect 317156 276350 317184 357750
rect 561508 313410 561536 674154
rect 579908 651137 579936 697983
rect 579894 651128 579950 651137
rect 579894 651063 579950 651072
rect 578790 627736 578846 627745
rect 578790 627671 578846 627680
rect 578804 627162 578832 627671
rect 578792 627156 578844 627162
rect 578792 627098 578844 627104
rect 579908 604217 579936 651063
rect 579894 604208 579950 604217
rect 579894 604143 579950 604152
rect 579158 580816 579214 580825
rect 579158 580751 579214 580760
rect 579172 334150 579200 580751
rect 579908 557297 579936 604143
rect 579894 557288 579950 557297
rect 579894 557223 579950 557232
rect 579250 533896 579306 533905
rect 579250 533831 579306 533840
rect 579264 358562 579292 533831
rect 579908 510377 579936 557223
rect 579894 510368 579950 510377
rect 579894 510303 579950 510312
rect 579342 486840 579398 486849
rect 579342 486775 579398 486784
rect 579252 358556 579304 358562
rect 579252 358498 579304 358504
rect 579356 358494 579384 486775
rect 579908 463457 579936 510303
rect 579894 463448 579950 463457
rect 579894 463383 579950 463392
rect 579434 439920 579490 439929
rect 579434 439855 579490 439864
rect 579344 358488 579396 358494
rect 579344 358430 579396 358436
rect 579448 354074 579476 439855
rect 579908 419506 579936 463383
rect 579724 419478 579936 419506
rect 579724 416537 579752 419478
rect 579710 416528 579766 416537
rect 579710 416463 579766 416472
rect 579724 409306 579752 416463
rect 579632 409278 579752 409306
rect 579526 393000 579582 393009
rect 579526 392935 579582 392944
rect 579436 354068 579488 354074
rect 579436 354010 579488 354016
rect 579160 334144 579212 334150
rect 579160 334086 579212 334092
rect 579540 313478 579568 392935
rect 579632 358426 579660 409278
rect 579620 358420 579672 358426
rect 579620 358362 579672 358368
rect 579528 313472 579580 313478
rect 579528 313414 579580 313420
rect 561496 313404 561548 313410
rect 561496 313346 561548 313352
rect 341800 276616 341852 276622
rect 341800 276558 341852 276564
rect 443090 276584 443146 276593
rect 326896 276548 326948 276554
rect 326896 276490 326948 276496
rect 337016 276548 337068 276554
rect 337016 276490 337068 276496
rect 317144 276344 317196 276350
rect 317144 276286 317196 276292
rect 326908 276282 326936 276490
rect 337028 276282 337056 276490
rect 316408 276276 316460 276282
rect 316408 276218 316460 276224
rect 326896 276276 326948 276282
rect 326896 276218 326948 276224
rect 337016 276276 337068 276282
rect 337016 276218 337068 276224
rect 316420 275942 316448 276218
rect 316408 275936 316460 275942
rect 316408 275878 316460 275884
rect 341812 273564 341840 276558
rect 347504 276548 347556 276554
rect 347504 276490 347556 276496
rect 357624 276548 357676 276554
rect 357624 276490 357676 276496
rect 365720 276548 365772 276554
rect 365720 276490 365772 276496
rect 403992 276548 404044 276554
rect 403992 276490 404044 276496
rect 419448 276548 419500 276554
rect 443090 276519 443092 276528
rect 419448 276490 419500 276496
rect 443144 276519 443146 276528
rect 453302 276584 453358 276593
rect 453302 276519 453358 276528
rect 443092 276490 443144 276496
rect 347516 276282 347544 276490
rect 357636 276282 357664 276490
rect 362776 276480 362828 276486
rect 362776 276422 362828 276428
rect 362788 276282 362816 276422
rect 347504 276276 347556 276282
rect 347504 276218 347556 276224
rect 357624 276276 357676 276282
rect 357624 276218 357676 276224
rect 362776 276276 362828 276282
rect 362776 276218 362828 276224
rect 365732 273564 365760 276490
rect 378232 276480 378284 276486
rect 378232 276422 378284 276428
rect 383384 276480 383436 276486
rect 383384 276422 383436 276428
rect 398840 276480 398892 276486
rect 398840 276422 398892 276428
rect 378244 276282 378272 276422
rect 383396 276282 383424 276422
rect 398852 276282 398880 276422
rect 404004 276282 404032 276490
rect 413928 276412 413980 276418
rect 413928 276354 413980 276360
rect 378232 276276 378284 276282
rect 378232 276218 378284 276224
rect 383384 276276 383436 276282
rect 383384 276218 383436 276224
rect 398840 276276 398892 276282
rect 398840 276218 398892 276224
rect 403992 276276 404044 276282
rect 403992 276218 404044 276224
rect 413940 273564 413968 276354
rect 419460 276282 419488 276490
rect 453316 276486 453344 276519
rect 429844 276480 429896 276486
rect 429844 276422 429896 276428
rect 435640 276480 435692 276486
rect 435732 276480 435784 276486
rect 435692 276428 435732 276434
rect 435640 276422 435784 276428
rect 453304 276480 453356 276486
rect 453304 276422 453356 276428
rect 454224 276480 454276 276486
rect 454224 276422 454276 276428
rect 429856 276282 429884 276422
rect 435652 276406 435772 276422
rect 438032 276344 438084 276350
rect 438032 276286 438084 276292
rect 419448 276276 419500 276282
rect 419448 276218 419500 276224
rect 429844 276276 429896 276282
rect 429844 276218 429896 276224
rect 438044 273564 438072 276286
rect 454236 276282 454264 276422
rect 454224 276276 454276 276282
rect 454224 276218 454276 276224
rect 461952 276276 462004 276282
rect 461952 276218 462004 276224
rect 461964 273564 461992 276218
rect 486056 276208 486108 276214
rect 486056 276150 486108 276156
rect 486068 273564 486096 276150
rect 510160 276140 510212 276146
rect 510160 276082 510212 276088
rect 510172 273564 510200 276082
rect 534264 276072 534316 276078
rect 534264 276014 534316 276020
rect 534276 273564 534304 276014
rect 558184 276004 558236 276010
rect 558184 275946 558236 275952
rect 558196 273564 558224 275946
rect 560852 272400 560904 272406
rect 560852 272342 560904 272348
rect 558644 272128 558696 272134
rect 558644 272070 558696 272076
rect 558656 267986 558684 272070
rect 558460 267980 558512 267986
rect 558460 267922 558512 267928
rect 558644 267980 558696 267986
rect 558644 267922 558696 267928
rect 558472 260522 558500 267922
rect 558472 260494 558592 260522
rect 558564 257582 558592 260494
rect 558552 257576 558604 257582
rect 558552 257518 558604 257524
rect 558644 257576 558696 257582
rect 558644 257518 558696 257524
rect 558656 250186 558684 257518
rect 558656 250158 558776 250186
rect 558748 247314 558776 250158
rect 558552 247308 558604 247314
rect 558552 247250 558604 247256
rect 558736 247308 558788 247314
rect 558736 247250 558788 247256
rect 558564 237046 558592 247250
rect 560864 237425 560892 272342
rect 560850 237416 560906 237425
rect 560850 237351 560906 237360
rect 558552 237040 558604 237046
rect 558552 236982 558604 236988
rect 558828 237040 558880 237046
rect 558828 236982 558880 236988
rect 558840 229770 558868 236982
rect 558828 229764 558880 229770
rect 558828 229706 558880 229712
rect 558736 229628 558788 229634
rect 558736 229570 558788 229576
rect 558748 219314 558776 229570
rect 558564 219286 558776 219314
rect 558564 209114 558592 219286
rect 558472 209086 558592 209114
rect 558472 203182 558500 209086
rect 558460 203176 558512 203182
rect 558460 203118 558512 203124
rect 558828 203176 558880 203182
rect 558828 203118 558880 203124
rect 558840 201929 558868 203118
rect 558826 201920 558882 201929
rect 558826 201855 558882 201864
rect 315670 163432 315726 163441
rect 315670 163367 315726 163376
rect 559378 130520 559434 130529
rect 559378 130455 559434 130464
rect 559392 125662 559420 130455
rect 558552 125656 558604 125662
rect 558552 125598 558604 125604
rect 559380 125656 559432 125662
rect 559380 125598 559432 125604
rect 315026 92440 315082 92449
rect 314200 92404 314252 92410
rect 315026 92375 315028 92384
rect 314200 92346 314252 92352
rect 315080 92375 315082 92384
rect 315028 92346 315080 92352
rect 314212 76022 314240 92346
rect 316500 81184 316552 81190
rect 316500 81126 316552 81132
rect 316512 76022 316540 81126
rect 558564 76022 558592 125598
rect 560850 95160 560906 95169
rect 560850 95095 560906 95104
rect 314200 76016 314252 76022
rect 314200 75958 314252 75964
rect 316500 76016 316552 76022
rect 316500 75958 316552 75964
rect 558552 76016 558604 76022
rect 558552 75958 558604 75964
rect 560864 75954 560892 95095
rect 560852 75948 560904 75954
rect 560852 75890 560904 75896
rect 314108 71868 314160 71874
rect 314108 71810 314160 71816
rect 313556 71800 313608 71806
rect 313556 71742 313608 71748
rect 331508 71534 331536 73644
rect 355612 71602 355640 73644
rect 379532 71670 379560 73644
rect 403636 71738 403664 73644
rect 427740 71874 427768 73644
rect 475948 72146 475976 73644
rect 475936 72140 475988 72146
rect 475936 72082 475988 72088
rect 499868 72010 499896 73644
rect 499856 72004 499908 72010
rect 499856 71946 499908 71952
rect 523972 71942 524000 73644
rect 548076 72078 548104 73644
rect 548064 72072 548116 72078
rect 548064 72014 548116 72020
rect 523960 71936 524012 71942
rect 523960 71878 524012 71884
rect 427728 71868 427780 71874
rect 427728 71810 427780 71816
rect 403624 71732 403676 71738
rect 403624 71674 403676 71680
rect 379520 71664 379572 71670
rect 379520 71606 379572 71612
rect 355600 71596 355652 71602
rect 355600 71538 355652 71544
rect 297272 71528 297324 71534
rect 297272 71470 297324 71476
rect 312360 71528 312412 71534
rect 312360 71470 312412 71476
rect 331496 71528 331548 71534
rect 331496 71470 331548 71476
rect 280160 71460 280212 71466
rect 280160 71402 280212 71408
rect 272432 71392 272484 71398
rect 272432 71334 272484 71340
rect 270592 3664 270644 3670
rect 270592 3606 270644 3612
rect 583392 3664 583444 3670
rect 583392 3606 583444 3612
rect 583404 480 583432 3606
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3606 667936 3662 667992
rect 2962 653540 3018 653576
rect 2962 653520 2964 653540
rect 2964 653520 3016 653540
rect 3016 653520 3018 653540
rect 2962 595992 3018 596048
rect 2962 538600 3018 538656
rect 2962 481072 3018 481128
rect 3698 610408 3754 610464
rect 257618 586064 257674 586120
rect 267738 586064 267794 586120
rect 3790 553016 3846 553072
rect 27250 581168 27306 581224
rect 24858 545536 24914 545592
rect 24950 509904 25006 509960
rect 3882 495488 3938 495544
rect 24858 473048 24914 473104
rect 24950 402056 25006 402112
rect 267922 386180 267924 386200
rect 267924 386180 267976 386200
rect 267976 386180 267978 386200
rect 267922 386144 267978 386180
rect 24766 199008 24822 199064
rect 24858 163376 24914 163432
rect 269302 547612 269304 547632
rect 269304 547612 269356 547632
rect 269356 547612 269358 547632
rect 269302 547576 269358 547612
rect 269302 511944 269358 512000
rect 269302 440680 269358 440736
rect 269302 405320 269358 405376
rect 270222 353776 270278 353832
rect 270038 348744 270094 348800
rect 269946 339904 270002 339960
rect 270130 339768 270186 339824
rect 269670 339632 269726 339688
rect 269854 335552 269910 335608
rect 270130 335552 270186 335608
rect 269394 329840 269450 329896
rect 175186 276684 175242 276720
rect 175186 276664 175188 276684
rect 175188 276664 175240 276684
rect 175240 276664 175242 276684
rect 185398 276664 185454 276720
rect 195794 276684 195850 276720
rect 195794 276664 195796 276684
rect 195796 276664 195848 276684
rect 195848 276664 195850 276684
rect 206006 276664 206062 276720
rect 216402 276684 216458 276720
rect 216402 276664 216404 276684
rect 216404 276664 216456 276684
rect 216456 276664 216458 276684
rect 226614 276664 226670 276720
rect 237010 276684 237066 276720
rect 237010 276664 237012 276684
rect 237012 276664 237064 276684
rect 237064 276664 237066 276684
rect 240046 276664 240102 276720
rect 26422 270272 26478 270328
rect 268382 237360 268438 237416
rect 26422 234640 26478 234696
rect 268382 201728 268438 201784
rect 269854 297336 269910 297392
rect 270406 345208 270462 345264
rect 270314 324400 270370 324456
rect 270314 297336 270370 297392
rect 270590 353776 270646 353832
rect 270590 350784 270646 350840
rect 270498 320728 270554 320784
rect 269854 236952 269910 237008
rect 270038 236952 270094 237008
rect 268566 166096 268622 166152
rect 270130 154536 270186 154592
rect 270406 154536 270462 154592
rect 270222 144236 270224 144256
rect 270224 144236 270276 144256
rect 270276 144236 270278 144256
rect 270222 144200 270278 144236
rect 270406 144200 270462 144256
rect 268290 130464 268346 130520
rect 24950 128016 25006 128072
rect 267922 95104 267978 95160
rect 24950 92384 25006 92440
rect 270682 333648 270738 333704
rect 270866 342624 270922 342680
rect 270774 317736 270830 317792
rect 272614 327528 272670 327584
rect 278134 386144 278190 386200
rect 298834 386436 298890 386472
rect 298834 386416 298836 386436
rect 298836 386416 298888 386436
rect 298888 386416 298890 386436
rect 309046 386416 309102 386472
rect 311530 352008 311586 352064
rect 312174 324944 312230 325000
rect 312082 318688 312138 318744
rect 312358 342896 312414 342952
rect 313554 339904 313610 339960
rect 313554 328208 313610 328264
rect 313554 327528 313610 327584
rect 313830 328208 313886 328264
rect 314014 345752 314070 345808
rect 314014 344528 314070 344584
rect 314014 333784 314070 333840
rect 314198 348744 314254 348800
rect 314198 344528 314254 344584
rect 314106 330928 314162 330984
rect 314382 402192 314438 402248
rect 314382 348744 314438 348800
rect 314290 336504 314346 336560
rect 579894 697992 579950 698048
rect 578514 674600 578570 674656
rect 463698 586492 463754 586528
rect 463698 586472 463700 586492
rect 463700 586472 463752 586492
rect 463752 586472 463754 586492
rect 473910 586472 473966 586528
rect 432786 586220 432842 586256
rect 432786 586200 432788 586220
rect 432788 586200 432840 586220
rect 432840 586200 432842 586220
rect 442906 586200 442962 586256
rect 315026 580660 315028 580680
rect 315028 580660 315080 580680
rect 315080 580660 315082 580680
rect 315026 580624 315082 580660
rect 315026 544892 315028 544912
rect 315028 544892 315080 544912
rect 315080 544892 315082 544912
rect 315026 544856 315082 544892
rect 560850 547712 560906 547768
rect 558918 512012 558974 512068
rect 315026 509668 315028 509688
rect 315028 509668 315080 509688
rect 315080 509668 315082 509688
rect 315026 509632 315082 509668
rect 315026 473048 315082 473104
rect 558918 440748 558974 440804
rect 560850 405320 560906 405376
rect 314474 321952 314530 322008
rect 315026 270272 315082 270328
rect 314290 234640 314346 234696
rect 315026 199008 315082 199064
rect 579894 651072 579950 651128
rect 578790 627680 578846 627736
rect 579894 604152 579950 604208
rect 579158 580760 579214 580816
rect 579894 557232 579950 557288
rect 579250 533840 579306 533896
rect 579894 510312 579950 510368
rect 579342 486784 579398 486840
rect 579894 463392 579950 463448
rect 579434 439864 579490 439920
rect 579710 416472 579766 416528
rect 579526 392944 579582 393000
rect 443090 276548 443146 276584
rect 443090 276528 443092 276548
rect 443092 276528 443144 276548
rect 443144 276528 443146 276548
rect 453302 276528 453358 276584
rect 560850 237360 560906 237416
rect 558826 201864 558882 201920
rect 315670 163376 315726 163432
rect 559378 130464 559434 130520
rect 315026 92404 315082 92440
rect 315026 92384 315028 92404
rect 315028 92384 315080 92404
rect 315080 92384 315082 92404
rect 560850 95104 560906 95160
<< metal3 >>
rect 579889 698050 579955 698053
rect 583520 698050 584960 698140
rect 579889 698048 584960 698050
rect 579889 697992 579894 698048
rect 579950 697992 584960 698048
rect 579889 697990 584960 697992
rect 579889 697987 579955 697990
rect 583520 697900 584960 697990
rect -960 696540 480 696780
rect 583520 686204 584960 686444
rect -960 682124 480 682364
rect 578509 674658 578575 674661
rect 583520 674658 584960 674748
rect 578509 674656 584960 674658
rect 578509 674600 578514 674656
rect 578570 674600 584960 674656
rect 578509 674598 584960 674600
rect 578509 674595 578575 674598
rect 583520 674508 584960 674598
rect -960 667994 480 668084
rect 3601 667994 3667 667997
rect -960 667992 3667 667994
rect -960 667936 3606 667992
rect 3662 667936 3667 667992
rect -960 667934 3667 667936
rect -960 667844 480 667934
rect 3601 667931 3667 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 2957 653578 3023 653581
rect -960 653576 3023 653578
rect -960 653520 2962 653576
rect 3018 653520 3023 653576
rect -960 653518 3023 653520
rect -960 653428 480 653518
rect 2957 653515 3023 653518
rect 579889 651130 579955 651133
rect 583520 651130 584960 651220
rect 579889 651128 584960 651130
rect 579889 651072 579894 651128
rect 579950 651072 584960 651128
rect 579889 651070 584960 651072
rect 579889 651067 579955 651070
rect 583520 650980 584960 651070
rect 583520 639284 584960 639524
rect -960 639012 480 639252
rect 578785 627738 578851 627741
rect 583520 627738 584960 627828
rect 578785 627736 584960 627738
rect 578785 627680 578790 627736
rect 578846 627680 584960 627736
rect 578785 627678 584960 627680
rect 578785 627675 578851 627678
rect 583520 627588 584960 627678
rect -960 624732 480 624972
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 3693 610466 3759 610469
rect -960 610464 3759 610466
rect -960 610408 3698 610464
rect 3754 610408 3759 610464
rect -960 610406 3759 610408
rect -960 610316 480 610406
rect 3693 610403 3759 610406
rect 579889 604210 579955 604213
rect 583520 604210 584960 604300
rect 579889 604208 584960 604210
rect 579889 604152 579894 604208
rect 579950 604152 584960 604208
rect 579889 604150 584960 604152
rect 579889 604147 579955 604150
rect 583520 604060 584960 604150
rect -960 596050 480 596140
rect 2957 596050 3023 596053
rect -960 596048 3023 596050
rect -960 595992 2962 596048
rect 3018 595992 3023 596048
rect -960 595990 3023 595992
rect -960 595900 480 595990
rect 2957 595987 3023 595990
rect 583520 592364 584960 592604
rect 463693 586530 463759 586533
rect 473905 586530 473971 586533
rect 463693 586528 473971 586530
rect 463693 586472 463698 586528
rect 463754 586472 473910 586528
rect 473966 586472 473971 586528
rect 463693 586470 473971 586472
rect 463693 586467 463759 586470
rect 473905 586467 473971 586470
rect 432781 586258 432847 586261
rect 442901 586258 442967 586261
rect 432781 586256 442967 586258
rect 432781 586200 432786 586256
rect 432842 586200 442906 586256
rect 442962 586200 442967 586256
rect 432781 586198 442967 586200
rect 432781 586195 432847 586198
rect 442901 586195 442967 586198
rect 257613 586122 257679 586125
rect 267733 586122 267799 586125
rect 257613 586120 267799 586122
rect 257613 586064 257618 586120
rect 257674 586064 267738 586120
rect 267794 586064 267799 586120
rect 257613 586062 267799 586064
rect 257613 586059 257679 586062
rect 267733 586059 267799 586062
rect -960 581620 480 581860
rect 27245 581226 27311 581229
rect 27245 581224 27354 581226
rect 27245 581168 27250 581224
rect 27306 581168 27354 581224
rect 27245 581163 27354 581168
rect 27294 580584 27354 581163
rect 579153 580818 579219 580821
rect 583520 580818 584960 580908
rect 579153 580816 584960 580818
rect 579153 580760 579158 580816
rect 579214 580760 584960 580816
rect 579153 580758 584960 580760
rect 579153 580755 579219 580758
rect 315021 580682 315087 580685
rect 315021 580680 318994 580682
rect 315021 580624 315026 580680
rect 315082 580624 318994 580680
rect 583520 580668 584960 580758
rect 315021 580622 318994 580624
rect 315021 580619 315087 580622
rect 318934 580584 318994 580622
rect 583520 568836 584960 569076
rect -960 567204 480 567444
rect 579889 557290 579955 557293
rect 583520 557290 584960 557380
rect 579889 557288 584960 557290
rect 579889 557232 579894 557288
rect 579950 557232 584960 557288
rect 579889 557230 584960 557232
rect 579889 557227 579955 557230
rect 583520 557140 584960 557230
rect -960 553074 480 553164
rect 3785 553074 3851 553077
rect -960 553072 3851 553074
rect -960 553016 3790 553072
rect 3846 553016 3851 553072
rect -960 553014 3851 553016
rect -960 552924 480 553014
rect 3785 553011 3851 553014
rect 560845 547770 560911 547773
rect 558870 547768 560911 547770
rect 558870 547712 560850 547768
rect 560906 547712 560911 547768
rect 558870 547710 560911 547712
rect 558870 547702 558930 547710
rect 560845 547707 560911 547710
rect 266524 547642 266922 547702
rect 558716 547642 558930 547702
rect 266862 547634 266922 547642
rect 269297 547634 269363 547637
rect 266862 547632 269363 547634
rect 266862 547576 269302 547632
rect 269358 547576 269363 547632
rect 266862 547574 269363 547576
rect 269297 547571 269363 547574
rect 24853 545594 24919 545597
rect 24853 545592 26802 545594
rect 24853 545536 24858 545592
rect 24914 545536 26802 545592
rect 24853 545534 26802 545536
rect 24853 545531 24919 545534
rect 26742 544952 26802 545534
rect 583520 545444 584960 545684
rect 315021 544914 315087 544917
rect 318934 544914 318994 544952
rect 315021 544912 318994 544914
rect 315021 544856 315026 544912
rect 315082 544856 318994 544912
rect 315021 544854 318994 544856
rect 315021 544851 315087 544854
rect -960 538658 480 538748
rect 2957 538658 3023 538661
rect -960 538656 3023 538658
rect -960 538600 2962 538656
rect 3018 538600 3023 538656
rect -960 538598 3023 538600
rect -960 538508 480 538598
rect 2957 538595 3023 538598
rect 579245 533898 579311 533901
rect 583520 533898 584960 533988
rect 579245 533896 584960 533898
rect 579245 533840 579250 533896
rect 579306 533840 584960 533896
rect 579245 533838 584960 533840
rect 579245 533835 579311 533838
rect 583520 533748 584960 533838
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 558913 512070 558979 512073
rect 266524 512010 267106 512070
rect 558716 512068 558979 512070
rect 558716 512012 558918 512068
rect 558974 512012 558979 512068
rect 558716 512010 558979 512012
rect 267046 512002 267106 512010
rect 558913 512007 558979 512010
rect 269297 512002 269363 512005
rect 267046 512000 269363 512002
rect 267046 511944 269302 512000
rect 269358 511944 269363 512000
rect 267046 511942 269363 511944
rect 269297 511939 269363 511942
rect 579889 510370 579955 510373
rect 583520 510370 584960 510460
rect 579889 510368 584960 510370
rect 579889 510312 579894 510368
rect 579950 510312 584960 510368
rect 579889 510310 584960 510312
rect 579889 510307 579955 510310
rect 583520 510220 584960 510310
rect -960 509812 480 510052
rect 24945 509962 25011 509965
rect 24945 509960 26802 509962
rect 24945 509904 24950 509960
rect 25006 509904 26802 509960
rect 24945 509902 26802 509904
rect 24945 509899 25011 509902
rect 26742 509320 26802 509902
rect 315021 509690 315087 509693
rect 315021 509688 318994 509690
rect 315021 509632 315026 509688
rect 315082 509632 318994 509688
rect 315021 509630 318994 509632
rect 315021 509627 315087 509630
rect 318934 509320 318994 509630
rect 583520 498524 584960 498764
rect -960 495546 480 495636
rect 3877 495546 3943 495549
rect -960 495544 3943 495546
rect -960 495488 3882 495544
rect 3938 495488 3943 495544
rect -960 495486 3943 495488
rect -960 495396 480 495486
rect 3877 495483 3943 495486
rect 579337 486842 579403 486845
rect 583520 486842 584960 486932
rect 579337 486840 584960 486842
rect 579337 486784 579342 486840
rect 579398 486784 584960 486840
rect 579337 486782 584960 486784
rect 579337 486779 579403 486782
rect 583520 486692 584960 486782
rect -960 481130 480 481220
rect 2957 481130 3023 481133
rect -960 481128 3023 481130
rect -960 481072 2962 481128
rect 3018 481072 3023 481128
rect -960 481070 3023 481072
rect -960 480980 480 481070
rect 2957 481067 3023 481070
rect 583520 474996 584960 475236
rect 24853 473106 24919 473109
rect 26742 473106 26802 473688
rect 24853 473104 26802 473106
rect 24853 473048 24858 473104
rect 24914 473048 26802 473104
rect 24853 473046 26802 473048
rect 315021 473106 315087 473109
rect 318934 473106 318994 473688
rect 315021 473104 318994 473106
rect 315021 473048 315026 473104
rect 315082 473048 318994 473104
rect 315021 473046 318994 473048
rect 24853 473043 24919 473046
rect 315021 473043 315087 473046
rect -960 466700 480 466940
rect 579889 463450 579955 463453
rect 583520 463450 584960 463540
rect 579889 463448 584960 463450
rect 579889 463392 579894 463448
rect 579950 463392 584960 463448
rect 579889 463390 584960 463392
rect 579889 463387 579955 463390
rect 583520 463300 584960 463390
rect -960 452284 480 452524
rect 583520 451604 584960 451844
rect 558913 440806 558979 440809
rect 266524 440746 266922 440806
rect 558716 440804 558979 440806
rect 558716 440748 558918 440804
rect 558974 440748 558979 440804
rect 558716 440746 558979 440748
rect 266862 440738 266922 440746
rect 558913 440743 558979 440746
rect 269297 440738 269363 440741
rect 266862 440736 269363 440738
rect 266862 440680 269302 440736
rect 269358 440680 269363 440736
rect 266862 440678 269363 440680
rect 269297 440675 269363 440678
rect 579429 439922 579495 439925
rect 583520 439922 584960 440012
rect 579429 439920 584960 439922
rect 579429 439864 579434 439920
rect 579490 439864 584960 439920
rect 579429 439862 584960 439864
rect 579429 439859 579495 439862
rect 583520 439772 584960 439862
rect -960 437868 480 438108
rect 583520 428076 584960 428316
rect -960 423588 480 423828
rect 579705 416530 579771 416533
rect 583520 416530 584960 416620
rect 579705 416528 584960 416530
rect 579705 416472 579710 416528
rect 579766 416472 584960 416528
rect 579705 416470 584960 416472
rect 579705 416467 579771 416470
rect 583520 416380 584960 416470
rect -960 409172 480 409412
rect 266524 405386 266922 405446
rect 558716 405386 559298 405446
rect 266862 405378 266922 405386
rect 269297 405378 269363 405381
rect 266862 405376 269363 405378
rect 266862 405320 269302 405376
rect 269358 405320 269363 405376
rect 266862 405318 269363 405320
rect 559238 405378 559298 405386
rect 560845 405378 560911 405381
rect 559238 405376 560911 405378
rect 559238 405320 560850 405376
rect 560906 405320 560911 405376
rect 559238 405318 560911 405320
rect 269297 405315 269363 405318
rect 560845 405315 560911 405318
rect 583520 404684 584960 404924
rect 24945 402114 25011 402117
rect 26742 402114 26802 402696
rect 314377 402250 314443 402253
rect 318934 402250 318994 402696
rect 314377 402248 318994 402250
rect 314377 402192 314382 402248
rect 314438 402192 318994 402248
rect 314377 402190 318994 402192
rect 314377 402187 314443 402190
rect 24945 402112 26802 402114
rect 24945 402056 24950 402112
rect 25006 402056 26802 402112
rect 24945 402054 26802 402056
rect 24945 402051 25011 402054
rect -960 394892 480 395132
rect 579521 393002 579587 393005
rect 583520 393002 584960 393092
rect 579521 393000 584960 393002
rect 579521 392944 579526 393000
rect 579582 392944 584960 393000
rect 579521 392942 584960 392944
rect 579521 392939 579587 392942
rect 583520 392852 584960 392942
rect 298829 386474 298895 386477
rect 309041 386474 309107 386477
rect 298829 386472 309107 386474
rect 298829 386416 298834 386472
rect 298890 386416 309046 386472
rect 309102 386416 309107 386472
rect 298829 386414 309107 386416
rect 298829 386411 298895 386414
rect 309041 386411 309107 386414
rect 267917 386202 267983 386205
rect 278129 386202 278195 386205
rect 267917 386200 278195 386202
rect 267917 386144 267922 386200
rect 267978 386144 278134 386200
rect 278190 386144 278195 386200
rect 267917 386142 278195 386144
rect 267917 386139 267983 386142
rect 278129 386139 278195 386142
rect 583520 381156 584960 381396
rect -960 380476 480 380716
rect 583520 369460 584960 369700
rect -960 366060 480 366300
rect 583520 357764 584960 358004
rect 270217 353834 270283 353837
rect 270585 353834 270651 353837
rect 272014 353834 272074 354348
rect 270217 353832 272074 353834
rect 270217 353776 270222 353832
rect 270278 353776 270590 353832
rect 270646 353776 272074 353832
rect 270217 353774 272074 353776
rect 270217 353771 270283 353774
rect 270585 353771 270651 353774
rect 311525 352066 311591 352069
rect 311525 352064 311634 352066
rect -960 351780 480 352020
rect 311525 352008 311530 352064
rect 311586 352008 311634 352064
rect 311525 352003 311634 352008
rect 311574 351628 311634 352003
rect 270585 350842 270651 350845
rect 272014 350842 272074 351356
rect 270585 350840 272074 350842
rect 270585 350784 270590 350840
rect 270646 350784 272074 350840
rect 270585 350782 272074 350784
rect 270585 350779 270651 350782
rect 270033 348802 270099 348805
rect 314193 348802 314259 348805
rect 314377 348802 314443 348805
rect 270033 348800 272074 348802
rect 270033 348744 270038 348800
rect 270094 348744 272074 348800
rect 270033 348742 272074 348744
rect 270033 348739 270099 348742
rect 272014 348364 272074 348742
rect 311942 348800 314443 348802
rect 311942 348744 314198 348800
rect 314254 348744 314382 348800
rect 314438 348744 314443 348800
rect 311942 348742 314443 348744
rect 311942 348636 312002 348742
rect 314193 348739 314259 348742
rect 314377 348739 314443 348742
rect 583520 345932 584960 346172
rect 314009 345810 314075 345813
rect 311942 345808 314075 345810
rect 311942 345752 314014 345808
rect 314070 345752 314075 345808
rect 311942 345750 314075 345752
rect 311942 345644 312002 345750
rect 314009 345747 314075 345750
rect 270401 345266 270467 345269
rect 272014 345266 272074 345372
rect 270401 345264 272074 345266
rect 270401 345208 270406 345264
rect 270462 345208 272074 345264
rect 270401 345206 272074 345208
rect 270401 345203 270467 345206
rect 314009 344586 314075 344589
rect 314193 344586 314259 344589
rect 314009 344584 314259 344586
rect 314009 344528 314014 344584
rect 314070 344528 314198 344584
rect 314254 344528 314259 344584
rect 314009 344526 314259 344528
rect 314009 344523 314075 344526
rect 314193 344523 314259 344526
rect 312353 342954 312419 342957
rect 311942 342952 312419 342954
rect 311942 342896 312358 342952
rect 312414 342896 312419 342952
rect 311942 342894 312419 342896
rect 270861 342682 270927 342685
rect 270861 342680 272074 342682
rect 270861 342624 270866 342680
rect 270922 342624 272074 342680
rect 311942 342652 312002 342894
rect 312353 342891 312419 342894
rect 270861 342622 272074 342624
rect 270861 342619 270927 342622
rect 272014 342108 272074 342622
rect 269941 339960 270007 339965
rect 313549 339962 313615 339965
rect 269941 339904 269946 339960
rect 270002 339904 270007 339960
rect 269941 339899 270007 339904
rect 311942 339960 313615 339962
rect 311942 339904 313554 339960
rect 313610 339904 313615 339960
rect 311942 339902 313615 339904
rect 269944 339826 270004 339899
rect 270125 339826 270191 339829
rect 269944 339824 270191 339826
rect 269944 339768 270130 339824
rect 270186 339768 270191 339824
rect 269944 339766 270191 339768
rect 270125 339763 270191 339766
rect 269665 339690 269731 339693
rect 269665 339688 272074 339690
rect 269665 339632 269670 339688
rect 269726 339632 272074 339688
rect 311942 339660 312002 339902
rect 313549 339899 313615 339902
rect 269665 339630 272074 339632
rect 269665 339627 269731 339630
rect 272014 339116 272074 339630
rect -960 337364 480 337604
rect 314285 336562 314351 336565
rect 311942 336560 314351 336562
rect 311942 336504 314290 336560
rect 314346 336504 314351 336560
rect 311942 336502 314351 336504
rect 311942 336396 312002 336502
rect 314285 336499 314351 336502
rect 269849 335610 269915 335613
rect 270125 335610 270191 335613
rect 272014 335610 272074 336124
rect 269849 335608 272074 335610
rect 269849 335552 269854 335608
rect 269910 335552 270130 335608
rect 270186 335552 272074 335608
rect 269849 335550 272074 335552
rect 269849 335547 269915 335550
rect 270125 335547 270191 335550
rect 583520 334236 584960 334476
rect 314009 333842 314075 333845
rect 311942 333840 314075 333842
rect 311942 333784 314014 333840
rect 314070 333784 314075 333840
rect 311942 333782 314075 333784
rect 270677 333706 270743 333709
rect 270677 333704 272074 333706
rect 270677 333648 270682 333704
rect 270738 333648 272074 333704
rect 270677 333646 272074 333648
rect 270677 333643 270743 333646
rect 272014 333132 272074 333646
rect 311942 333404 312002 333782
rect 314009 333779 314075 333782
rect 314101 330986 314167 330989
rect 311942 330984 314167 330986
rect 311942 330928 314106 330984
rect 314162 330928 314167 330984
rect 311942 330926 314167 330928
rect 311942 330412 312002 330926
rect 314101 330923 314167 330926
rect 269389 329898 269455 329901
rect 272014 329898 272074 330140
rect 269389 329896 272074 329898
rect 269389 329840 269394 329896
rect 269450 329840 272074 329896
rect 269389 329838 272074 329840
rect 269389 329835 269455 329838
rect 313549 328266 313615 328269
rect 313825 328266 313891 328269
rect 313549 328264 313891 328266
rect 313549 328208 313554 328264
rect 313610 328208 313830 328264
rect 313886 328208 313891 328264
rect 313549 328206 313891 328208
rect 313549 328203 313615 328206
rect 313825 328203 313891 328206
rect 272609 327586 272675 327589
rect 313549 327586 313615 327589
rect 272566 327584 272675 327586
rect 272566 327528 272614 327584
rect 272670 327528 272675 327584
rect 272566 327523 272675 327528
rect 311942 327584 313615 327586
rect 311942 327528 313554 327584
rect 313610 327528 313615 327584
rect 311942 327526 313615 327528
rect 272566 327148 272626 327523
rect 311942 327420 312002 327526
rect 313549 327523 313615 327526
rect 312169 325002 312235 325005
rect 311942 325000 312235 325002
rect 311942 324944 312174 325000
rect 312230 324944 312235 325000
rect 311942 324942 312235 324944
rect 270309 324458 270375 324461
rect 270309 324456 272074 324458
rect 270309 324400 270314 324456
rect 270370 324400 272074 324456
rect 311942 324428 312002 324942
rect 312169 324939 312235 324942
rect 270309 324398 272074 324400
rect 270309 324395 270375 324398
rect 272014 323884 272074 324398
rect -960 322948 480 323188
rect 583520 322540 584960 322780
rect 314469 322010 314535 322013
rect 311942 322008 314535 322010
rect 311942 321952 314474 322008
rect 314530 321952 314535 322008
rect 311942 321950 314535 321952
rect 311942 321436 312002 321950
rect 314469 321947 314535 321950
rect 270493 320786 270559 320789
rect 272014 320786 272074 320892
rect 270493 320784 272074 320786
rect 270493 320728 270498 320784
rect 270554 320728 272074 320784
rect 270493 320726 272074 320728
rect 270493 320723 270559 320726
rect 312077 318746 312143 318749
rect 311942 318744 312143 318746
rect 311942 318688 312082 318744
rect 312138 318688 312143 318744
rect 311942 318686 312143 318688
rect 311942 318172 312002 318686
rect 312077 318683 312143 318686
rect 270769 317794 270835 317797
rect 272014 317794 272074 317900
rect 270769 317792 272074 317794
rect 270769 317736 270774 317792
rect 270830 317736 272074 317792
rect 270769 317734 272074 317736
rect 270769 317731 270835 317734
rect 583520 310708 584960 310948
rect -960 308668 480 308908
rect 583520 299012 584960 299252
rect 269849 297394 269915 297397
rect 270309 297394 270375 297397
rect 269849 297392 270375 297394
rect 269849 297336 269854 297392
rect 269910 297336 270314 297392
rect 270370 297336 270375 297392
rect 269849 297334 270375 297336
rect 269849 297331 269915 297334
rect 270309 297331 270375 297334
rect -960 294252 480 294492
rect 583520 287316 584960 287556
rect -960 279972 480 280212
rect 175181 276722 175247 276725
rect 185393 276722 185459 276725
rect 175181 276720 185459 276722
rect 175181 276664 175186 276720
rect 175242 276664 185398 276720
rect 185454 276664 185459 276720
rect 175181 276662 185459 276664
rect 175181 276659 175247 276662
rect 185393 276659 185459 276662
rect 195789 276722 195855 276725
rect 206001 276722 206067 276725
rect 195789 276720 206067 276722
rect 195789 276664 195794 276720
rect 195850 276664 206006 276720
rect 206062 276664 206067 276720
rect 195789 276662 206067 276664
rect 195789 276659 195855 276662
rect 206001 276659 206067 276662
rect 216397 276722 216463 276725
rect 226609 276722 226675 276725
rect 216397 276720 226675 276722
rect 216397 276664 216402 276720
rect 216458 276664 226614 276720
rect 226670 276664 226675 276720
rect 216397 276662 226675 276664
rect 216397 276659 216463 276662
rect 226609 276659 226675 276662
rect 237005 276722 237071 276725
rect 240041 276722 240107 276725
rect 237005 276720 240107 276722
rect 237005 276664 237010 276720
rect 237066 276664 240046 276720
rect 240102 276664 240107 276720
rect 237005 276662 240107 276664
rect 237005 276659 237071 276662
rect 240041 276659 240107 276662
rect 443085 276586 443151 276589
rect 453297 276586 453363 276589
rect 443085 276584 453363 276586
rect 443085 276528 443090 276584
rect 443146 276528 453302 276584
rect 453358 276528 453363 276584
rect 443085 276526 453363 276528
rect 443085 276523 443151 276526
rect 453297 276523 453363 276526
rect 583520 275620 584960 275860
rect 26417 270330 26483 270333
rect 315021 270330 315087 270333
rect 26417 270328 26772 270330
rect 26417 270272 26422 270328
rect 26478 270272 26772 270328
rect 26417 270270 26772 270272
rect 315021 270328 318964 270330
rect 315021 270272 315026 270328
rect 315082 270272 318964 270328
rect 315021 270270 318964 270272
rect 26417 270267 26483 270270
rect 315021 270267 315087 270270
rect -960 265556 480 265796
rect 583520 263788 584960 264028
rect 583520 252092 584960 252332
rect -960 251140 480 251380
rect 583520 240396 584960 240636
rect 268377 237418 268443 237421
rect 560845 237418 560911 237421
rect 266524 237416 268443 237418
rect 266524 237360 268382 237416
rect 268438 237360 268443 237416
rect 266524 237358 268443 237360
rect 558716 237416 560911 237418
rect 558716 237360 560850 237416
rect 560906 237360 560911 237416
rect 558716 237358 560911 237360
rect 268377 237355 268443 237358
rect 560845 237355 560911 237358
rect -960 236860 480 237100
rect 269849 237010 269915 237013
rect 270033 237010 270099 237013
rect 269849 237008 270099 237010
rect 269849 236952 269854 237008
rect 269910 236952 270038 237008
rect 270094 236952 270099 237008
rect 269849 236950 270099 236952
rect 269849 236947 269915 236950
rect 270033 236947 270099 236950
rect 26417 234698 26483 234701
rect 314285 234698 314351 234701
rect 26417 234696 26772 234698
rect 26417 234640 26422 234696
rect 26478 234640 26772 234696
rect 26417 234638 26772 234640
rect 314285 234696 318964 234698
rect 314285 234640 314290 234696
rect 314346 234640 318964 234696
rect 314285 234638 318964 234640
rect 26417 234635 26483 234638
rect 314285 234635 314351 234638
rect 583520 228700 584960 228940
rect -960 222444 480 222684
rect 583520 216868 584960 217108
rect -960 208028 480 208268
rect 583520 205172 584960 205412
rect 558821 201922 558887 201925
rect 558821 201920 558930 201922
rect 558821 201864 558826 201920
rect 558882 201864 558930 201920
rect 558821 201859 558930 201864
rect 268377 201786 268443 201789
rect 558870 201786 558930 201859
rect 266524 201784 268443 201786
rect 266524 201728 268382 201784
rect 268438 201728 268443 201784
rect 266524 201726 268443 201728
rect 558716 201726 558930 201786
rect 268377 201723 268443 201726
rect 24761 199066 24827 199069
rect 315021 199066 315087 199069
rect 24761 199064 26772 199066
rect 24761 199008 24766 199064
rect 24822 199008 26772 199064
rect 24761 199006 26772 199008
rect 315021 199064 318964 199066
rect 315021 199008 315026 199064
rect 315082 199008 318964 199064
rect 315021 199006 318964 199008
rect 24761 199003 24827 199006
rect 315021 199003 315087 199006
rect -960 193748 480 193988
rect 583520 193476 584960 193716
rect 583520 181780 584960 182020
rect -960 179332 480 179572
rect 583520 169948 584960 170188
rect 268561 166154 268627 166157
rect 266524 166152 268627 166154
rect 266524 166096 268566 166152
rect 268622 166096 268627 166152
rect 266524 166094 268627 166096
rect 268561 166091 268627 166094
rect -960 164916 480 165156
rect 24853 163434 24919 163437
rect 315665 163434 315731 163437
rect 24853 163432 26772 163434
rect 24853 163376 24858 163432
rect 24914 163376 26772 163432
rect 24853 163374 26772 163376
rect 315665 163432 318964 163434
rect 315665 163376 315670 163432
rect 315726 163376 318964 163432
rect 315665 163374 318964 163376
rect 24853 163371 24919 163374
rect 315665 163371 315731 163374
rect 583520 158252 584960 158492
rect 270125 154594 270191 154597
rect 270401 154594 270467 154597
rect 270125 154592 270467 154594
rect 270125 154536 270130 154592
rect 270186 154536 270406 154592
rect 270462 154536 270467 154592
rect 270125 154534 270467 154536
rect 270125 154531 270191 154534
rect 270401 154531 270467 154534
rect -960 150636 480 150876
rect 583520 146556 584960 146796
rect 270217 144258 270283 144261
rect 270401 144258 270467 144261
rect 270217 144256 270467 144258
rect 270217 144200 270222 144256
rect 270278 144200 270406 144256
rect 270462 144200 270467 144256
rect 270217 144198 270467 144200
rect 270217 144195 270283 144198
rect 270401 144195 270467 144198
rect -960 136220 480 136460
rect 583520 134724 584960 134964
rect 268285 130522 268351 130525
rect 559373 130522 559439 130525
rect 266524 130520 268351 130522
rect 266524 130464 268290 130520
rect 268346 130464 268351 130520
rect 266524 130462 268351 130464
rect 558716 130520 559439 130522
rect 558716 130464 559378 130520
rect 559434 130464 559439 130520
rect 558716 130462 559439 130464
rect 268285 130459 268351 130462
rect 559373 130459 559439 130462
rect 24945 128074 25011 128077
rect 24945 128072 26772 128074
rect 24945 128016 24950 128072
rect 25006 128016 26772 128072
rect 24945 128014 26772 128016
rect 24945 128011 25011 128014
rect 583520 123028 584960 123268
rect -960 121940 480 122180
rect 583520 111332 584960 111572
rect -960 107524 480 107764
rect 583520 99636 584960 99876
rect 267917 95162 267983 95165
rect 560845 95162 560911 95165
rect 266524 95160 267983 95162
rect 266524 95104 267922 95160
rect 267978 95104 267983 95160
rect 266524 95102 267983 95104
rect 558716 95160 560911 95162
rect 558716 95104 560850 95160
rect 560906 95104 560911 95160
rect 558716 95102 560911 95104
rect 267917 95099 267983 95102
rect 560845 95099 560911 95102
rect -960 93108 480 93348
rect 24945 92442 25011 92445
rect 315021 92442 315087 92445
rect 24945 92440 26772 92442
rect 24945 92384 24950 92440
rect 25006 92384 26772 92440
rect 24945 92382 26772 92384
rect 315021 92440 318964 92442
rect 315021 92384 315026 92440
rect 315082 92384 318964 92440
rect 315021 92382 318964 92384
rect 24945 92379 25011 92382
rect 315021 92379 315087 92382
rect 583520 87804 584960 88044
rect -960 78828 480 79068
rect 583520 76108 584960 76348
rect -960 64412 480 64652
rect 583520 64412 584960 64652
rect 583520 52716 584960 52956
rect -960 49996 480 50236
rect 583520 40884 584960 41124
rect -960 35716 480 35956
rect 583520 29188 584960 29428
rect -960 21300 480 21540
rect 583520 17492 584960 17732
rect -960 7020 480 7260
rect 583520 5796 584960 6036
<< metal4 >>
rect -8576 711418 -7976 711440
rect -8576 711182 -8394 711418
rect -8158 711182 -7976 711418
rect -8576 711098 -7976 711182
rect -8576 710862 -8394 711098
rect -8158 710862 -7976 711098
rect -8576 -6926 -7976 710862
rect 591900 711418 592500 711440
rect 591900 711182 592082 711418
rect 592318 711182 592500 711418
rect 591900 711098 592500 711182
rect 591900 710862 592082 711098
rect 592318 710862 592500 711098
rect -7636 710478 -7036 710500
rect -7636 710242 -7454 710478
rect -7218 710242 -7036 710478
rect -7636 710158 -7036 710242
rect -7636 709922 -7454 710158
rect -7218 709922 -7036 710158
rect -7636 -5986 -7036 709922
rect 590960 710478 591560 710500
rect 590960 710242 591142 710478
rect 591378 710242 591560 710478
rect 590960 710158 591560 710242
rect 590960 709922 591142 710158
rect 591378 709922 591560 710158
rect -6696 709538 -6096 709560
rect -6696 709302 -6514 709538
rect -6278 709302 -6096 709538
rect -6696 709218 -6096 709302
rect -6696 708982 -6514 709218
rect -6278 708982 -6096 709218
rect -6696 -5046 -6096 708982
rect 590020 709538 590620 709560
rect 590020 709302 590202 709538
rect 590438 709302 590620 709538
rect 590020 709218 590620 709302
rect 590020 708982 590202 709218
rect 590438 708982 590620 709218
rect -5756 708598 -5156 708620
rect -5756 708362 -5574 708598
rect -5338 708362 -5156 708598
rect -5756 708278 -5156 708362
rect -5756 708042 -5574 708278
rect -5338 708042 -5156 708278
rect -5756 -4106 -5156 708042
rect 589080 708598 589680 708620
rect 589080 708362 589262 708598
rect 589498 708362 589680 708598
rect 589080 708278 589680 708362
rect 589080 708042 589262 708278
rect 589498 708042 589680 708278
rect -4816 707658 -4216 707680
rect -4816 707422 -4634 707658
rect -4398 707422 -4216 707658
rect -4816 707338 -4216 707422
rect -4816 707102 -4634 707338
rect -4398 707102 -4216 707338
rect -4816 -3166 -4216 707102
rect 588140 707658 588740 707680
rect 588140 707422 588322 707658
rect 588558 707422 588740 707658
rect 588140 707338 588740 707422
rect 588140 707102 588322 707338
rect 588558 707102 588740 707338
rect -3876 706718 -3276 706740
rect -3876 706482 -3694 706718
rect -3458 706482 -3276 706718
rect -3876 706398 -3276 706482
rect -3876 706162 -3694 706398
rect -3458 706162 -3276 706398
rect -3876 -2226 -3276 706162
rect 587200 706718 587800 706740
rect 587200 706482 587382 706718
rect 587618 706482 587800 706718
rect 587200 706398 587800 706482
rect 587200 706162 587382 706398
rect 587618 706162 587800 706398
rect -2936 705778 -2336 705800
rect -2936 705542 -2754 705778
rect -2518 705542 -2336 705778
rect -2936 705458 -2336 705542
rect -2936 705222 -2754 705458
rect -2518 705222 -2336 705458
rect -2936 668454 -2336 705222
rect -2936 668218 -2754 668454
rect -2518 668218 -2336 668454
rect -2936 668134 -2336 668218
rect -2936 667898 -2754 668134
rect -2518 667898 -2336 668134
rect -2936 632454 -2336 667898
rect -2936 632218 -2754 632454
rect -2518 632218 -2336 632454
rect -2936 632134 -2336 632218
rect -2936 631898 -2754 632134
rect -2518 631898 -2336 632134
rect -2936 596454 -2336 631898
rect -2936 596218 -2754 596454
rect -2518 596218 -2336 596454
rect -2936 596134 -2336 596218
rect -2936 595898 -2754 596134
rect -2518 595898 -2336 596134
rect -2936 560454 -2336 595898
rect -2936 560218 -2754 560454
rect -2518 560218 -2336 560454
rect -2936 560134 -2336 560218
rect -2936 559898 -2754 560134
rect -2518 559898 -2336 560134
rect -2936 524454 -2336 559898
rect -2936 524218 -2754 524454
rect -2518 524218 -2336 524454
rect -2936 524134 -2336 524218
rect -2936 523898 -2754 524134
rect -2518 523898 -2336 524134
rect -2936 488454 -2336 523898
rect -2936 488218 -2754 488454
rect -2518 488218 -2336 488454
rect -2936 488134 -2336 488218
rect -2936 487898 -2754 488134
rect -2518 487898 -2336 488134
rect -2936 452454 -2336 487898
rect -2936 452218 -2754 452454
rect -2518 452218 -2336 452454
rect -2936 452134 -2336 452218
rect -2936 451898 -2754 452134
rect -2518 451898 -2336 452134
rect -2936 416454 -2336 451898
rect -2936 416218 -2754 416454
rect -2518 416218 -2336 416454
rect -2936 416134 -2336 416218
rect -2936 415898 -2754 416134
rect -2518 415898 -2336 416134
rect -2936 380454 -2336 415898
rect -2936 380218 -2754 380454
rect -2518 380218 -2336 380454
rect -2936 380134 -2336 380218
rect -2936 379898 -2754 380134
rect -2518 379898 -2336 380134
rect -2936 344454 -2336 379898
rect -2936 344218 -2754 344454
rect -2518 344218 -2336 344454
rect -2936 344134 -2336 344218
rect -2936 343898 -2754 344134
rect -2518 343898 -2336 344134
rect -2936 308454 -2336 343898
rect -2936 308218 -2754 308454
rect -2518 308218 -2336 308454
rect -2936 308134 -2336 308218
rect -2936 307898 -2754 308134
rect -2518 307898 -2336 308134
rect -2936 272454 -2336 307898
rect -2936 272218 -2754 272454
rect -2518 272218 -2336 272454
rect -2936 272134 -2336 272218
rect -2936 271898 -2754 272134
rect -2518 271898 -2336 272134
rect -2936 236454 -2336 271898
rect -2936 236218 -2754 236454
rect -2518 236218 -2336 236454
rect -2936 236134 -2336 236218
rect -2936 235898 -2754 236134
rect -2518 235898 -2336 236134
rect -2936 200454 -2336 235898
rect -2936 200218 -2754 200454
rect -2518 200218 -2336 200454
rect -2936 200134 -2336 200218
rect -2936 199898 -2754 200134
rect -2518 199898 -2336 200134
rect -2936 164454 -2336 199898
rect -2936 164218 -2754 164454
rect -2518 164218 -2336 164454
rect -2936 164134 -2336 164218
rect -2936 163898 -2754 164134
rect -2518 163898 -2336 164134
rect -2936 128454 -2336 163898
rect -2936 128218 -2754 128454
rect -2518 128218 -2336 128454
rect -2936 128134 -2336 128218
rect -2936 127898 -2754 128134
rect -2518 127898 -2336 128134
rect -2936 92454 -2336 127898
rect -2936 92218 -2754 92454
rect -2518 92218 -2336 92454
rect -2936 92134 -2336 92218
rect -2936 91898 -2754 92134
rect -2518 91898 -2336 92134
rect -2936 56454 -2336 91898
rect -2936 56218 -2754 56454
rect -2518 56218 -2336 56454
rect -2936 56134 -2336 56218
rect -2936 55898 -2754 56134
rect -2518 55898 -2336 56134
rect -2936 20454 -2336 55898
rect -2936 20218 -2754 20454
rect -2518 20218 -2336 20454
rect -2936 20134 -2336 20218
rect -2936 19898 -2754 20134
rect -2518 19898 -2336 20134
rect -2936 -1286 -2336 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705800
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2936 -1522 -2754 -1286
rect -2518 -1522 -2336 -1286
rect -2936 -1606 -2336 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 -2336 -1606
rect -2936 -1864 -2336 -1842
rect 804 -1864 1404 -902
rect 18804 705778 19404 705800
rect 18804 705542 18986 705778
rect 19222 705542 19404 705778
rect 18804 705458 19404 705542
rect 18804 705222 18986 705458
rect 19222 705222 19404 705458
rect 18804 668454 19404 705222
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 36804 704838 37404 705800
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 584916 37404 613898
rect 54804 705778 55404 705800
rect 54804 705542 54986 705778
rect 55222 705542 55404 705778
rect 54804 705458 55404 705542
rect 54804 705222 54986 705458
rect 55222 705222 55404 705458
rect 54804 668454 55404 705222
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 584916 55404 595898
rect 72804 704838 73404 705800
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 614454 73404 649898
rect 72804 614218 72986 614454
rect 73222 614218 73404 614454
rect 72804 614134 73404 614218
rect 72804 613898 72986 614134
rect 73222 613898 73404 614134
rect 72804 584916 73404 613898
rect 90804 705778 91404 705800
rect 90804 705542 90986 705778
rect 91222 705542 91404 705778
rect 90804 705458 91404 705542
rect 90804 705222 90986 705458
rect 91222 705222 91404 705458
rect 90804 668454 91404 705222
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 632454 91404 667898
rect 90804 632218 90986 632454
rect 91222 632218 91404 632454
rect 90804 632134 91404 632218
rect 90804 631898 90986 632134
rect 91222 631898 91404 632134
rect 90804 596454 91404 631898
rect 90804 596218 90986 596454
rect 91222 596218 91404 596454
rect 90804 596134 91404 596218
rect 90804 595898 90986 596134
rect 91222 595898 91404 596134
rect 90804 584916 91404 595898
rect 108804 704838 109404 705800
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 650454 109404 685898
rect 108804 650218 108986 650454
rect 109222 650218 109404 650454
rect 108804 650134 109404 650218
rect 108804 649898 108986 650134
rect 109222 649898 109404 650134
rect 108804 614454 109404 649898
rect 108804 614218 108986 614454
rect 109222 614218 109404 614454
rect 108804 614134 109404 614218
rect 108804 613898 108986 614134
rect 109222 613898 109404 614134
rect 108804 584916 109404 613898
rect 126804 705778 127404 705800
rect 126804 705542 126986 705778
rect 127222 705542 127404 705778
rect 126804 705458 127404 705542
rect 126804 705222 126986 705458
rect 127222 705222 127404 705458
rect 126804 668454 127404 705222
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 632454 127404 667898
rect 126804 632218 126986 632454
rect 127222 632218 127404 632454
rect 126804 632134 127404 632218
rect 126804 631898 126986 632134
rect 127222 631898 127404 632134
rect 126804 596454 127404 631898
rect 126804 596218 126986 596454
rect 127222 596218 127404 596454
rect 126804 596134 127404 596218
rect 126804 595898 126986 596134
rect 127222 595898 127404 596134
rect 126804 584916 127404 595898
rect 144804 704838 145404 705800
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 144804 584916 145404 613898
rect 162804 705778 163404 705800
rect 162804 705542 162986 705778
rect 163222 705542 163404 705778
rect 162804 705458 163404 705542
rect 162804 705222 162986 705458
rect 163222 705222 163404 705458
rect 162804 668454 163404 705222
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 162804 584916 163404 595898
rect 180804 704838 181404 705800
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 584916 181404 613898
rect 198804 705778 199404 705800
rect 198804 705542 198986 705778
rect 199222 705542 199404 705778
rect 198804 705458 199404 705542
rect 198804 705222 198986 705458
rect 199222 705222 199404 705458
rect 198804 668454 199404 705222
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 632454 199404 667898
rect 198804 632218 198986 632454
rect 199222 632218 199404 632454
rect 198804 632134 199404 632218
rect 198804 631898 198986 632134
rect 199222 631898 199404 632134
rect 198804 596454 199404 631898
rect 198804 596218 198986 596454
rect 199222 596218 199404 596454
rect 198804 596134 199404 596218
rect 198804 595898 198986 596134
rect 199222 595898 199404 596134
rect 198804 584916 199404 595898
rect 216804 704838 217404 705800
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 650454 217404 685898
rect 216804 650218 216986 650454
rect 217222 650218 217404 650454
rect 216804 650134 217404 650218
rect 216804 649898 216986 650134
rect 217222 649898 217404 650134
rect 216804 614454 217404 649898
rect 216804 614218 216986 614454
rect 217222 614218 217404 614454
rect 216804 614134 217404 614218
rect 216804 613898 216986 614134
rect 217222 613898 217404 614134
rect 216804 584916 217404 613898
rect 234804 705778 235404 705800
rect 234804 705542 234986 705778
rect 235222 705542 235404 705778
rect 234804 705458 235404 705542
rect 234804 705222 234986 705458
rect 235222 705222 235404 705458
rect 234804 668454 235404 705222
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 632454 235404 667898
rect 234804 632218 234986 632454
rect 235222 632218 235404 632454
rect 234804 632134 235404 632218
rect 234804 631898 234986 632134
rect 235222 631898 235404 632134
rect 234804 596454 235404 631898
rect 234804 596218 234986 596454
rect 235222 596218 235404 596454
rect 234804 596134 235404 596218
rect 234804 595898 234986 596134
rect 235222 595898 235404 596134
rect 234804 584916 235404 595898
rect 252804 704838 253404 705800
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 650454 253404 685898
rect 252804 650218 252986 650454
rect 253222 650218 253404 650454
rect 252804 650134 253404 650218
rect 252804 649898 252986 650134
rect 253222 649898 253404 650134
rect 252804 614454 253404 649898
rect 252804 614218 252986 614454
rect 253222 614218 253404 614454
rect 252804 614134 253404 614218
rect 252804 613898 252986 614134
rect 253222 613898 253404 614134
rect 252804 584916 253404 613898
rect 270804 705778 271404 705800
rect 270804 705542 270986 705778
rect 271222 705542 271404 705778
rect 270804 705458 271404 705542
rect 270804 705222 270986 705458
rect 271222 705222 271404 705458
rect 270804 668454 271404 705222
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 270804 596454 271404 631898
rect 270804 596218 270986 596454
rect 271222 596218 271404 596454
rect 270804 596134 271404 596218
rect 270804 595898 270986 596134
rect 271222 595898 271404 596134
rect 47088 578454 47408 578476
rect 47088 578218 47130 578454
rect 47366 578218 47408 578454
rect 47088 578134 47408 578218
rect 47088 577898 47130 578134
rect 47366 577898 47408 578134
rect 47088 577876 47408 577898
rect 77808 578454 78128 578476
rect 77808 578218 77850 578454
rect 78086 578218 78128 578454
rect 77808 578134 78128 578218
rect 77808 577898 77850 578134
rect 78086 577898 78128 578134
rect 77808 577876 78128 577898
rect 108528 578454 108848 578476
rect 108528 578218 108570 578454
rect 108806 578218 108848 578454
rect 108528 578134 108848 578218
rect 108528 577898 108570 578134
rect 108806 577898 108848 578134
rect 108528 577876 108848 577898
rect 139248 578454 139568 578476
rect 139248 578218 139290 578454
rect 139526 578218 139568 578454
rect 139248 578134 139568 578218
rect 139248 577898 139290 578134
rect 139526 577898 139568 578134
rect 139248 577876 139568 577898
rect 169968 578454 170288 578476
rect 169968 578218 170010 578454
rect 170246 578218 170288 578454
rect 169968 578134 170288 578218
rect 169968 577898 170010 578134
rect 170246 577898 170288 578134
rect 169968 577876 170288 577898
rect 200688 578454 201008 578476
rect 200688 578218 200730 578454
rect 200966 578218 201008 578454
rect 200688 578134 201008 578218
rect 200688 577898 200730 578134
rect 200966 577898 201008 578134
rect 200688 577876 201008 577898
rect 231408 578454 231728 578476
rect 231408 578218 231450 578454
rect 231686 578218 231728 578454
rect 231408 578134 231728 578218
rect 231408 577898 231450 578134
rect 231686 577898 231728 578134
rect 231408 577876 231728 577898
rect 262128 578454 262448 578476
rect 262128 578218 262170 578454
rect 262406 578218 262448 578454
rect 262128 578134 262448 578218
rect 262128 577898 262170 578134
rect 262406 577898 262448 578134
rect 262128 577876 262448 577898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 31728 560454 32048 560476
rect 31728 560218 31770 560454
rect 32006 560218 32048 560454
rect 31728 560134 32048 560218
rect 31728 559898 31770 560134
rect 32006 559898 32048 560134
rect 31728 559876 32048 559898
rect 62448 560454 62768 560476
rect 62448 560218 62490 560454
rect 62726 560218 62768 560454
rect 62448 560134 62768 560218
rect 62448 559898 62490 560134
rect 62726 559898 62768 560134
rect 62448 559876 62768 559898
rect 93168 560454 93488 560476
rect 93168 560218 93210 560454
rect 93446 560218 93488 560454
rect 93168 560134 93488 560218
rect 93168 559898 93210 560134
rect 93446 559898 93488 560134
rect 93168 559876 93488 559898
rect 123888 560454 124208 560476
rect 123888 560218 123930 560454
rect 124166 560218 124208 560454
rect 123888 560134 124208 560218
rect 123888 559898 123930 560134
rect 124166 559898 124208 560134
rect 123888 559876 124208 559898
rect 154608 560454 154928 560476
rect 154608 560218 154650 560454
rect 154886 560218 154928 560454
rect 154608 560134 154928 560218
rect 154608 559898 154650 560134
rect 154886 559898 154928 560134
rect 154608 559876 154928 559898
rect 185328 560454 185648 560476
rect 185328 560218 185370 560454
rect 185606 560218 185648 560454
rect 185328 560134 185648 560218
rect 185328 559898 185370 560134
rect 185606 559898 185648 560134
rect 185328 559876 185648 559898
rect 216048 560454 216368 560476
rect 216048 560218 216090 560454
rect 216326 560218 216368 560454
rect 216048 560134 216368 560218
rect 216048 559898 216090 560134
rect 216326 559898 216368 560134
rect 216048 559876 216368 559898
rect 246768 560454 247088 560476
rect 246768 560218 246810 560454
rect 247046 560218 247088 560454
rect 246768 560134 247088 560218
rect 246768 559898 246810 560134
rect 247046 559898 247088 560134
rect 246768 559876 247088 559898
rect 270804 560454 271404 595898
rect 270804 560218 270986 560454
rect 271222 560218 271404 560454
rect 270804 560134 271404 560218
rect 270804 559898 270986 560134
rect 271222 559898 271404 560134
rect 47088 542454 47408 542476
rect 47088 542218 47130 542454
rect 47366 542218 47408 542454
rect 47088 542134 47408 542218
rect 47088 541898 47130 542134
rect 47366 541898 47408 542134
rect 47088 541876 47408 541898
rect 77808 542454 78128 542476
rect 77808 542218 77850 542454
rect 78086 542218 78128 542454
rect 77808 542134 78128 542218
rect 77808 541898 77850 542134
rect 78086 541898 78128 542134
rect 77808 541876 78128 541898
rect 108528 542454 108848 542476
rect 108528 542218 108570 542454
rect 108806 542218 108848 542454
rect 108528 542134 108848 542218
rect 108528 541898 108570 542134
rect 108806 541898 108848 542134
rect 108528 541876 108848 541898
rect 139248 542454 139568 542476
rect 139248 542218 139290 542454
rect 139526 542218 139568 542454
rect 139248 542134 139568 542218
rect 139248 541898 139290 542134
rect 139526 541898 139568 542134
rect 139248 541876 139568 541898
rect 169968 542454 170288 542476
rect 169968 542218 170010 542454
rect 170246 542218 170288 542454
rect 169968 542134 170288 542218
rect 169968 541898 170010 542134
rect 170246 541898 170288 542134
rect 169968 541876 170288 541898
rect 200688 542454 201008 542476
rect 200688 542218 200730 542454
rect 200966 542218 201008 542454
rect 200688 542134 201008 542218
rect 200688 541898 200730 542134
rect 200966 541898 201008 542134
rect 200688 541876 201008 541898
rect 231408 542454 231728 542476
rect 231408 542218 231450 542454
rect 231686 542218 231728 542454
rect 231408 542134 231728 542218
rect 231408 541898 231450 542134
rect 231686 541898 231728 542134
rect 231408 541876 231728 541898
rect 262128 542454 262448 542476
rect 262128 542218 262170 542454
rect 262406 542218 262448 542454
rect 262128 542134 262448 542218
rect 262128 541898 262170 542134
rect 262406 541898 262448 542134
rect 262128 541876 262448 541898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 31728 524454 32048 524476
rect 31728 524218 31770 524454
rect 32006 524218 32048 524454
rect 31728 524134 32048 524218
rect 31728 523898 31770 524134
rect 32006 523898 32048 524134
rect 31728 523876 32048 523898
rect 62448 524454 62768 524476
rect 62448 524218 62490 524454
rect 62726 524218 62768 524454
rect 62448 524134 62768 524218
rect 62448 523898 62490 524134
rect 62726 523898 62768 524134
rect 62448 523876 62768 523898
rect 93168 524454 93488 524476
rect 93168 524218 93210 524454
rect 93446 524218 93488 524454
rect 93168 524134 93488 524218
rect 93168 523898 93210 524134
rect 93446 523898 93488 524134
rect 93168 523876 93488 523898
rect 123888 524454 124208 524476
rect 123888 524218 123930 524454
rect 124166 524218 124208 524454
rect 123888 524134 124208 524218
rect 123888 523898 123930 524134
rect 124166 523898 124208 524134
rect 123888 523876 124208 523898
rect 154608 524454 154928 524476
rect 154608 524218 154650 524454
rect 154886 524218 154928 524454
rect 154608 524134 154928 524218
rect 154608 523898 154650 524134
rect 154886 523898 154928 524134
rect 154608 523876 154928 523898
rect 185328 524454 185648 524476
rect 185328 524218 185370 524454
rect 185606 524218 185648 524454
rect 185328 524134 185648 524218
rect 185328 523898 185370 524134
rect 185606 523898 185648 524134
rect 185328 523876 185648 523898
rect 216048 524454 216368 524476
rect 216048 524218 216090 524454
rect 216326 524218 216368 524454
rect 216048 524134 216368 524218
rect 216048 523898 216090 524134
rect 216326 523898 216368 524134
rect 216048 523876 216368 523898
rect 246768 524454 247088 524476
rect 246768 524218 246810 524454
rect 247046 524218 247088 524454
rect 246768 524134 247088 524218
rect 246768 523898 246810 524134
rect 247046 523898 247088 524134
rect 246768 523876 247088 523898
rect 270804 524454 271404 559898
rect 270804 524218 270986 524454
rect 271222 524218 271404 524454
rect 270804 524134 271404 524218
rect 270804 523898 270986 524134
rect 271222 523898 271404 524134
rect 47088 506454 47408 506476
rect 47088 506218 47130 506454
rect 47366 506218 47408 506454
rect 47088 506134 47408 506218
rect 47088 505898 47130 506134
rect 47366 505898 47408 506134
rect 47088 505876 47408 505898
rect 77808 506454 78128 506476
rect 77808 506218 77850 506454
rect 78086 506218 78128 506454
rect 77808 506134 78128 506218
rect 77808 505898 77850 506134
rect 78086 505898 78128 506134
rect 77808 505876 78128 505898
rect 108528 506454 108848 506476
rect 108528 506218 108570 506454
rect 108806 506218 108848 506454
rect 108528 506134 108848 506218
rect 108528 505898 108570 506134
rect 108806 505898 108848 506134
rect 108528 505876 108848 505898
rect 139248 506454 139568 506476
rect 139248 506218 139290 506454
rect 139526 506218 139568 506454
rect 139248 506134 139568 506218
rect 139248 505898 139290 506134
rect 139526 505898 139568 506134
rect 139248 505876 139568 505898
rect 169968 506454 170288 506476
rect 169968 506218 170010 506454
rect 170246 506218 170288 506454
rect 169968 506134 170288 506218
rect 169968 505898 170010 506134
rect 170246 505898 170288 506134
rect 169968 505876 170288 505898
rect 200688 506454 201008 506476
rect 200688 506218 200730 506454
rect 200966 506218 201008 506454
rect 200688 506134 201008 506218
rect 200688 505898 200730 506134
rect 200966 505898 201008 506134
rect 200688 505876 201008 505898
rect 231408 506454 231728 506476
rect 231408 506218 231450 506454
rect 231686 506218 231728 506454
rect 231408 506134 231728 506218
rect 231408 505898 231450 506134
rect 231686 505898 231728 506134
rect 231408 505876 231728 505898
rect 262128 506454 262448 506476
rect 262128 506218 262170 506454
rect 262406 506218 262448 506454
rect 262128 506134 262448 506218
rect 262128 505898 262170 506134
rect 262406 505898 262448 506134
rect 262128 505876 262448 505898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 31728 488454 32048 488476
rect 31728 488218 31770 488454
rect 32006 488218 32048 488454
rect 31728 488134 32048 488218
rect 31728 487898 31770 488134
rect 32006 487898 32048 488134
rect 31728 487876 32048 487898
rect 62448 488454 62768 488476
rect 62448 488218 62490 488454
rect 62726 488218 62768 488454
rect 62448 488134 62768 488218
rect 62448 487898 62490 488134
rect 62726 487898 62768 488134
rect 62448 487876 62768 487898
rect 93168 488454 93488 488476
rect 93168 488218 93210 488454
rect 93446 488218 93488 488454
rect 93168 488134 93488 488218
rect 93168 487898 93210 488134
rect 93446 487898 93488 488134
rect 93168 487876 93488 487898
rect 123888 488454 124208 488476
rect 123888 488218 123930 488454
rect 124166 488218 124208 488454
rect 123888 488134 124208 488218
rect 123888 487898 123930 488134
rect 124166 487898 124208 488134
rect 123888 487876 124208 487898
rect 154608 488454 154928 488476
rect 154608 488218 154650 488454
rect 154886 488218 154928 488454
rect 154608 488134 154928 488218
rect 154608 487898 154650 488134
rect 154886 487898 154928 488134
rect 154608 487876 154928 487898
rect 185328 488454 185648 488476
rect 185328 488218 185370 488454
rect 185606 488218 185648 488454
rect 185328 488134 185648 488218
rect 185328 487898 185370 488134
rect 185606 487898 185648 488134
rect 185328 487876 185648 487898
rect 216048 488454 216368 488476
rect 216048 488218 216090 488454
rect 216326 488218 216368 488454
rect 216048 488134 216368 488218
rect 216048 487898 216090 488134
rect 216326 487898 216368 488134
rect 216048 487876 216368 487898
rect 246768 488454 247088 488476
rect 246768 488218 246810 488454
rect 247046 488218 247088 488454
rect 246768 488134 247088 488218
rect 246768 487898 246810 488134
rect 247046 487898 247088 488134
rect 246768 487876 247088 487898
rect 270804 488454 271404 523898
rect 270804 488218 270986 488454
rect 271222 488218 271404 488454
rect 270804 488134 271404 488218
rect 270804 487898 270986 488134
rect 271222 487898 271404 488134
rect 47088 470454 47408 470476
rect 47088 470218 47130 470454
rect 47366 470218 47408 470454
rect 47088 470134 47408 470218
rect 47088 469898 47130 470134
rect 47366 469898 47408 470134
rect 47088 469876 47408 469898
rect 77808 470454 78128 470476
rect 77808 470218 77850 470454
rect 78086 470218 78128 470454
rect 77808 470134 78128 470218
rect 77808 469898 77850 470134
rect 78086 469898 78128 470134
rect 77808 469876 78128 469898
rect 108528 470454 108848 470476
rect 108528 470218 108570 470454
rect 108806 470218 108848 470454
rect 108528 470134 108848 470218
rect 108528 469898 108570 470134
rect 108806 469898 108848 470134
rect 108528 469876 108848 469898
rect 139248 470454 139568 470476
rect 139248 470218 139290 470454
rect 139526 470218 139568 470454
rect 139248 470134 139568 470218
rect 139248 469898 139290 470134
rect 139526 469898 139568 470134
rect 139248 469876 139568 469898
rect 169968 470454 170288 470476
rect 169968 470218 170010 470454
rect 170246 470218 170288 470454
rect 169968 470134 170288 470218
rect 169968 469898 170010 470134
rect 170246 469898 170288 470134
rect 169968 469876 170288 469898
rect 200688 470454 201008 470476
rect 200688 470218 200730 470454
rect 200966 470218 201008 470454
rect 200688 470134 201008 470218
rect 200688 469898 200730 470134
rect 200966 469898 201008 470134
rect 200688 469876 201008 469898
rect 231408 470454 231728 470476
rect 231408 470218 231450 470454
rect 231686 470218 231728 470454
rect 231408 470134 231728 470218
rect 231408 469898 231450 470134
rect 231686 469898 231728 470134
rect 231408 469876 231728 469898
rect 262128 470454 262448 470476
rect 262128 470218 262170 470454
rect 262406 470218 262448 470454
rect 262128 470134 262448 470218
rect 262128 469898 262170 470134
rect 262406 469898 262448 470134
rect 262128 469876 262448 469898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 31728 452454 32048 452476
rect 31728 452218 31770 452454
rect 32006 452218 32048 452454
rect 31728 452134 32048 452218
rect 31728 451898 31770 452134
rect 32006 451898 32048 452134
rect 31728 451876 32048 451898
rect 62448 452454 62768 452476
rect 62448 452218 62490 452454
rect 62726 452218 62768 452454
rect 62448 452134 62768 452218
rect 62448 451898 62490 452134
rect 62726 451898 62768 452134
rect 62448 451876 62768 451898
rect 93168 452454 93488 452476
rect 93168 452218 93210 452454
rect 93446 452218 93488 452454
rect 93168 452134 93488 452218
rect 93168 451898 93210 452134
rect 93446 451898 93488 452134
rect 93168 451876 93488 451898
rect 123888 452454 124208 452476
rect 123888 452218 123930 452454
rect 124166 452218 124208 452454
rect 123888 452134 124208 452218
rect 123888 451898 123930 452134
rect 124166 451898 124208 452134
rect 123888 451876 124208 451898
rect 154608 452454 154928 452476
rect 154608 452218 154650 452454
rect 154886 452218 154928 452454
rect 154608 452134 154928 452218
rect 154608 451898 154650 452134
rect 154886 451898 154928 452134
rect 154608 451876 154928 451898
rect 185328 452454 185648 452476
rect 185328 452218 185370 452454
rect 185606 452218 185648 452454
rect 185328 452134 185648 452218
rect 185328 451898 185370 452134
rect 185606 451898 185648 452134
rect 185328 451876 185648 451898
rect 216048 452454 216368 452476
rect 216048 452218 216090 452454
rect 216326 452218 216368 452454
rect 216048 452134 216368 452218
rect 216048 451898 216090 452134
rect 216326 451898 216368 452134
rect 216048 451876 216368 451898
rect 246768 452454 247088 452476
rect 246768 452218 246810 452454
rect 247046 452218 247088 452454
rect 246768 452134 247088 452218
rect 246768 451898 246810 452134
rect 247046 451898 247088 452134
rect 246768 451876 247088 451898
rect 270804 452454 271404 487898
rect 270804 452218 270986 452454
rect 271222 452218 271404 452454
rect 270804 452134 271404 452218
rect 270804 451898 270986 452134
rect 271222 451898 271404 452134
rect 47088 434454 47408 434476
rect 47088 434218 47130 434454
rect 47366 434218 47408 434454
rect 47088 434134 47408 434218
rect 47088 433898 47130 434134
rect 47366 433898 47408 434134
rect 47088 433876 47408 433898
rect 77808 434454 78128 434476
rect 77808 434218 77850 434454
rect 78086 434218 78128 434454
rect 77808 434134 78128 434218
rect 77808 433898 77850 434134
rect 78086 433898 78128 434134
rect 77808 433876 78128 433898
rect 108528 434454 108848 434476
rect 108528 434218 108570 434454
rect 108806 434218 108848 434454
rect 108528 434134 108848 434218
rect 108528 433898 108570 434134
rect 108806 433898 108848 434134
rect 108528 433876 108848 433898
rect 139248 434454 139568 434476
rect 139248 434218 139290 434454
rect 139526 434218 139568 434454
rect 139248 434134 139568 434218
rect 139248 433898 139290 434134
rect 139526 433898 139568 434134
rect 139248 433876 139568 433898
rect 169968 434454 170288 434476
rect 169968 434218 170010 434454
rect 170246 434218 170288 434454
rect 169968 434134 170288 434218
rect 169968 433898 170010 434134
rect 170246 433898 170288 434134
rect 169968 433876 170288 433898
rect 200688 434454 201008 434476
rect 200688 434218 200730 434454
rect 200966 434218 201008 434454
rect 200688 434134 201008 434218
rect 200688 433898 200730 434134
rect 200966 433898 201008 434134
rect 200688 433876 201008 433898
rect 231408 434454 231728 434476
rect 231408 434218 231450 434454
rect 231686 434218 231728 434454
rect 231408 434134 231728 434218
rect 231408 433898 231450 434134
rect 231686 433898 231728 434134
rect 231408 433876 231728 433898
rect 262128 434454 262448 434476
rect 262128 434218 262170 434454
rect 262406 434218 262448 434454
rect 262128 434134 262448 434218
rect 262128 433898 262170 434134
rect 262406 433898 262448 434134
rect 262128 433876 262448 433898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 31728 416454 32048 416476
rect 31728 416218 31770 416454
rect 32006 416218 32048 416454
rect 31728 416134 32048 416218
rect 31728 415898 31770 416134
rect 32006 415898 32048 416134
rect 31728 415876 32048 415898
rect 62448 416454 62768 416476
rect 62448 416218 62490 416454
rect 62726 416218 62768 416454
rect 62448 416134 62768 416218
rect 62448 415898 62490 416134
rect 62726 415898 62768 416134
rect 62448 415876 62768 415898
rect 93168 416454 93488 416476
rect 93168 416218 93210 416454
rect 93446 416218 93488 416454
rect 93168 416134 93488 416218
rect 93168 415898 93210 416134
rect 93446 415898 93488 416134
rect 93168 415876 93488 415898
rect 123888 416454 124208 416476
rect 123888 416218 123930 416454
rect 124166 416218 124208 416454
rect 123888 416134 124208 416218
rect 123888 415898 123930 416134
rect 124166 415898 124208 416134
rect 123888 415876 124208 415898
rect 154608 416454 154928 416476
rect 154608 416218 154650 416454
rect 154886 416218 154928 416454
rect 154608 416134 154928 416218
rect 154608 415898 154650 416134
rect 154886 415898 154928 416134
rect 154608 415876 154928 415898
rect 185328 416454 185648 416476
rect 185328 416218 185370 416454
rect 185606 416218 185648 416454
rect 185328 416134 185648 416218
rect 185328 415898 185370 416134
rect 185606 415898 185648 416134
rect 185328 415876 185648 415898
rect 216048 416454 216368 416476
rect 216048 416218 216090 416454
rect 216326 416218 216368 416454
rect 216048 416134 216368 416218
rect 216048 415898 216090 416134
rect 216326 415898 216368 416134
rect 216048 415876 216368 415898
rect 246768 416454 247088 416476
rect 246768 416218 246810 416454
rect 247046 416218 247088 416454
rect 246768 416134 247088 416218
rect 246768 415898 246810 416134
rect 247046 415898 247088 416134
rect 246768 415876 247088 415898
rect 270804 416454 271404 451898
rect 270804 416218 270986 416454
rect 271222 416218 271404 416454
rect 270804 416134 271404 416218
rect 270804 415898 270986 416134
rect 271222 415898 271404 416134
rect 47088 398454 47408 398476
rect 47088 398218 47130 398454
rect 47366 398218 47408 398454
rect 47088 398134 47408 398218
rect 47088 397898 47130 398134
rect 47366 397898 47408 398134
rect 47088 397876 47408 397898
rect 77808 398454 78128 398476
rect 77808 398218 77850 398454
rect 78086 398218 78128 398454
rect 77808 398134 78128 398218
rect 77808 397898 77850 398134
rect 78086 397898 78128 398134
rect 77808 397876 78128 397898
rect 108528 398454 108848 398476
rect 108528 398218 108570 398454
rect 108806 398218 108848 398454
rect 108528 398134 108848 398218
rect 108528 397898 108570 398134
rect 108806 397898 108848 398134
rect 108528 397876 108848 397898
rect 139248 398454 139568 398476
rect 139248 398218 139290 398454
rect 139526 398218 139568 398454
rect 139248 398134 139568 398218
rect 139248 397898 139290 398134
rect 139526 397898 139568 398134
rect 139248 397876 139568 397898
rect 169968 398454 170288 398476
rect 169968 398218 170010 398454
rect 170246 398218 170288 398454
rect 169968 398134 170288 398218
rect 169968 397898 170010 398134
rect 170246 397898 170288 398134
rect 169968 397876 170288 397898
rect 200688 398454 201008 398476
rect 200688 398218 200730 398454
rect 200966 398218 201008 398454
rect 200688 398134 201008 398218
rect 200688 397898 200730 398134
rect 200966 397898 201008 398134
rect 200688 397876 201008 397898
rect 231408 398454 231728 398476
rect 231408 398218 231450 398454
rect 231686 398218 231728 398454
rect 231408 398134 231728 398218
rect 231408 397898 231450 398134
rect 231686 397898 231728 398134
rect 231408 397876 231728 397898
rect 262128 398454 262448 398476
rect 262128 398218 262170 398454
rect 262406 398218 262448 398454
rect 262128 398134 262448 398218
rect 262128 397898 262170 398134
rect 262406 397898 262448 398134
rect 262128 397876 262448 397898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 36804 362454 37404 382916
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 274600 37404 289898
rect 54804 380454 55404 382916
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 274600 55404 307898
rect 72804 362454 73404 382916
rect 72804 362218 72986 362454
rect 73222 362218 73404 362454
rect 72804 362134 73404 362218
rect 72804 361898 72986 362134
rect 73222 361898 73404 362134
rect 72804 326454 73404 361898
rect 72804 326218 72986 326454
rect 73222 326218 73404 326454
rect 72804 326134 73404 326218
rect 72804 325898 72986 326134
rect 73222 325898 73404 326134
rect 72804 290454 73404 325898
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 274600 73404 289898
rect 90804 380454 91404 382916
rect 90804 380218 90986 380454
rect 91222 380218 91404 380454
rect 90804 380134 91404 380218
rect 90804 379898 90986 380134
rect 91222 379898 91404 380134
rect 90804 344454 91404 379898
rect 90804 344218 90986 344454
rect 91222 344218 91404 344454
rect 90804 344134 91404 344218
rect 90804 343898 90986 344134
rect 91222 343898 91404 344134
rect 90804 308454 91404 343898
rect 90804 308218 90986 308454
rect 91222 308218 91404 308454
rect 90804 308134 91404 308218
rect 90804 307898 90986 308134
rect 91222 307898 91404 308134
rect 90804 274600 91404 307898
rect 108804 362454 109404 382916
rect 108804 362218 108986 362454
rect 109222 362218 109404 362454
rect 108804 362134 109404 362218
rect 108804 361898 108986 362134
rect 109222 361898 109404 362134
rect 108804 326454 109404 361898
rect 108804 326218 108986 326454
rect 109222 326218 109404 326454
rect 108804 326134 109404 326218
rect 108804 325898 108986 326134
rect 109222 325898 109404 326134
rect 108804 290454 109404 325898
rect 108804 290218 108986 290454
rect 109222 290218 109404 290454
rect 108804 290134 109404 290218
rect 108804 289898 108986 290134
rect 109222 289898 109404 290134
rect 108804 274600 109404 289898
rect 126804 380454 127404 382916
rect 126804 380218 126986 380454
rect 127222 380218 127404 380454
rect 126804 380134 127404 380218
rect 126804 379898 126986 380134
rect 127222 379898 127404 380134
rect 126804 344454 127404 379898
rect 126804 344218 126986 344454
rect 127222 344218 127404 344454
rect 126804 344134 127404 344218
rect 126804 343898 126986 344134
rect 127222 343898 127404 344134
rect 126804 308454 127404 343898
rect 126804 308218 126986 308454
rect 127222 308218 127404 308454
rect 126804 308134 127404 308218
rect 126804 307898 126986 308134
rect 127222 307898 127404 308134
rect 126804 274600 127404 307898
rect 144804 362454 145404 382916
rect 144804 362218 144986 362454
rect 145222 362218 145404 362454
rect 144804 362134 145404 362218
rect 144804 361898 144986 362134
rect 145222 361898 145404 362134
rect 144804 326454 145404 361898
rect 144804 326218 144986 326454
rect 145222 326218 145404 326454
rect 144804 326134 145404 326218
rect 144804 325898 144986 326134
rect 145222 325898 145404 326134
rect 144804 290454 145404 325898
rect 144804 290218 144986 290454
rect 145222 290218 145404 290454
rect 144804 290134 145404 290218
rect 144804 289898 144986 290134
rect 145222 289898 145404 290134
rect 144804 274600 145404 289898
rect 162804 380454 163404 382916
rect 162804 380218 162986 380454
rect 163222 380218 163404 380454
rect 162804 380134 163404 380218
rect 162804 379898 162986 380134
rect 163222 379898 163404 380134
rect 162804 344454 163404 379898
rect 162804 344218 162986 344454
rect 163222 344218 163404 344454
rect 162804 344134 163404 344218
rect 162804 343898 162986 344134
rect 163222 343898 163404 344134
rect 162804 308454 163404 343898
rect 162804 308218 162986 308454
rect 163222 308218 163404 308454
rect 162804 308134 163404 308218
rect 162804 307898 162986 308134
rect 163222 307898 163404 308134
rect 162804 274600 163404 307898
rect 180804 362454 181404 382916
rect 180804 362218 180986 362454
rect 181222 362218 181404 362454
rect 180804 362134 181404 362218
rect 180804 361898 180986 362134
rect 181222 361898 181404 362134
rect 180804 326454 181404 361898
rect 180804 326218 180986 326454
rect 181222 326218 181404 326454
rect 180804 326134 181404 326218
rect 180804 325898 180986 326134
rect 181222 325898 181404 326134
rect 180804 290454 181404 325898
rect 180804 290218 180986 290454
rect 181222 290218 181404 290454
rect 180804 290134 181404 290218
rect 180804 289898 180986 290134
rect 181222 289898 181404 290134
rect 180804 274600 181404 289898
rect 198804 380454 199404 382916
rect 198804 380218 198986 380454
rect 199222 380218 199404 380454
rect 198804 380134 199404 380218
rect 198804 379898 198986 380134
rect 199222 379898 199404 380134
rect 198804 344454 199404 379898
rect 198804 344218 198986 344454
rect 199222 344218 199404 344454
rect 198804 344134 199404 344218
rect 198804 343898 198986 344134
rect 199222 343898 199404 344134
rect 198804 308454 199404 343898
rect 198804 308218 198986 308454
rect 199222 308218 199404 308454
rect 198804 308134 199404 308218
rect 198804 307898 198986 308134
rect 199222 307898 199404 308134
rect 198804 274600 199404 307898
rect 216804 362454 217404 382916
rect 216804 362218 216986 362454
rect 217222 362218 217404 362454
rect 216804 362134 217404 362218
rect 216804 361898 216986 362134
rect 217222 361898 217404 362134
rect 216804 326454 217404 361898
rect 216804 326218 216986 326454
rect 217222 326218 217404 326454
rect 216804 326134 217404 326218
rect 216804 325898 216986 326134
rect 217222 325898 217404 326134
rect 216804 290454 217404 325898
rect 216804 290218 216986 290454
rect 217222 290218 217404 290454
rect 216804 290134 217404 290218
rect 216804 289898 216986 290134
rect 217222 289898 217404 290134
rect 216804 274600 217404 289898
rect 234804 380454 235404 382916
rect 234804 380218 234986 380454
rect 235222 380218 235404 380454
rect 234804 380134 235404 380218
rect 234804 379898 234986 380134
rect 235222 379898 235404 380134
rect 234804 344454 235404 379898
rect 234804 344218 234986 344454
rect 235222 344218 235404 344454
rect 234804 344134 235404 344218
rect 234804 343898 234986 344134
rect 235222 343898 235404 344134
rect 234804 308454 235404 343898
rect 234804 308218 234986 308454
rect 235222 308218 235404 308454
rect 234804 308134 235404 308218
rect 234804 307898 234986 308134
rect 235222 307898 235404 308134
rect 234804 274600 235404 307898
rect 252804 362454 253404 382916
rect 252804 362218 252986 362454
rect 253222 362218 253404 362454
rect 252804 362134 253404 362218
rect 252804 361898 252986 362134
rect 253222 361898 253404 362134
rect 252804 326454 253404 361898
rect 270804 380454 271404 415898
rect 270804 380218 270986 380454
rect 271222 380218 271404 380454
rect 270804 380134 271404 380218
rect 270804 379898 270986 380134
rect 271222 379898 271404 380134
rect 270804 356560 271404 379898
rect 288804 704838 289404 705800
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 578454 289404 613898
rect 288804 578218 288986 578454
rect 289222 578218 289404 578454
rect 288804 578134 289404 578218
rect 288804 577898 288986 578134
rect 289222 577898 289404 578134
rect 288804 542454 289404 577898
rect 288804 542218 288986 542454
rect 289222 542218 289404 542454
rect 288804 542134 289404 542218
rect 288804 541898 288986 542134
rect 289222 541898 289404 542134
rect 288804 506454 289404 541898
rect 288804 506218 288986 506454
rect 289222 506218 289404 506454
rect 288804 506134 289404 506218
rect 288804 505898 288986 506134
rect 289222 505898 289404 506134
rect 288804 470454 289404 505898
rect 288804 470218 288986 470454
rect 289222 470218 289404 470454
rect 288804 470134 289404 470218
rect 288804 469898 288986 470134
rect 289222 469898 289404 470134
rect 288804 434454 289404 469898
rect 288804 434218 288986 434454
rect 289222 434218 289404 434454
rect 288804 434134 289404 434218
rect 288804 433898 288986 434134
rect 289222 433898 289404 434134
rect 288804 398454 289404 433898
rect 288804 398218 288986 398454
rect 289222 398218 289404 398454
rect 288804 398134 289404 398218
rect 288804 397898 288986 398134
rect 289222 397898 289404 398134
rect 288804 362454 289404 397898
rect 288804 362218 288986 362454
rect 289222 362218 289404 362454
rect 288804 362134 289404 362218
rect 288804 361898 288986 362134
rect 289222 361898 289404 362134
rect 288804 356560 289404 361898
rect 306804 705778 307404 705800
rect 306804 705542 306986 705778
rect 307222 705542 307404 705778
rect 306804 705458 307404 705542
rect 306804 705222 306986 705458
rect 307222 705222 307404 705458
rect 306804 668454 307404 705222
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 632454 307404 667898
rect 306804 632218 306986 632454
rect 307222 632218 307404 632454
rect 306804 632134 307404 632218
rect 306804 631898 306986 632134
rect 307222 631898 307404 632134
rect 306804 596454 307404 631898
rect 306804 596218 306986 596454
rect 307222 596218 307404 596454
rect 306804 596134 307404 596218
rect 306804 595898 306986 596134
rect 307222 595898 307404 596134
rect 306804 560454 307404 595898
rect 324804 704838 325404 705800
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 650454 325404 685898
rect 324804 650218 324986 650454
rect 325222 650218 325404 650454
rect 324804 650134 325404 650218
rect 324804 649898 324986 650134
rect 325222 649898 325404 650134
rect 324804 614454 325404 649898
rect 324804 614218 324986 614454
rect 325222 614218 325404 614454
rect 324804 614134 325404 614218
rect 324804 613898 324986 614134
rect 325222 613898 325404 614134
rect 324804 584916 325404 613898
rect 342804 705778 343404 705800
rect 342804 705542 342986 705778
rect 343222 705542 343404 705778
rect 342804 705458 343404 705542
rect 342804 705222 342986 705458
rect 343222 705222 343404 705458
rect 342804 668454 343404 705222
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 632454 343404 667898
rect 342804 632218 342986 632454
rect 343222 632218 343404 632454
rect 342804 632134 343404 632218
rect 342804 631898 342986 632134
rect 343222 631898 343404 632134
rect 342804 596454 343404 631898
rect 342804 596218 342986 596454
rect 343222 596218 343404 596454
rect 342804 596134 343404 596218
rect 342804 595898 342986 596134
rect 343222 595898 343404 596134
rect 342804 584916 343404 595898
rect 360804 704838 361404 705800
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 650454 361404 685898
rect 360804 650218 360986 650454
rect 361222 650218 361404 650454
rect 360804 650134 361404 650218
rect 360804 649898 360986 650134
rect 361222 649898 361404 650134
rect 360804 614454 361404 649898
rect 360804 614218 360986 614454
rect 361222 614218 361404 614454
rect 360804 614134 361404 614218
rect 360804 613898 360986 614134
rect 361222 613898 361404 614134
rect 360804 584916 361404 613898
rect 378804 705778 379404 705800
rect 378804 705542 378986 705778
rect 379222 705542 379404 705778
rect 378804 705458 379404 705542
rect 378804 705222 378986 705458
rect 379222 705222 379404 705458
rect 378804 668454 379404 705222
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 632454 379404 667898
rect 378804 632218 378986 632454
rect 379222 632218 379404 632454
rect 378804 632134 379404 632218
rect 378804 631898 378986 632134
rect 379222 631898 379404 632134
rect 378804 596454 379404 631898
rect 378804 596218 378986 596454
rect 379222 596218 379404 596454
rect 378804 596134 379404 596218
rect 378804 595898 378986 596134
rect 379222 595898 379404 596134
rect 378804 584916 379404 595898
rect 396804 704838 397404 705800
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 396804 614454 397404 649898
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 396804 584916 397404 613898
rect 414804 705778 415404 705800
rect 414804 705542 414986 705778
rect 415222 705542 415404 705778
rect 414804 705458 415404 705542
rect 414804 705222 414986 705458
rect 415222 705222 415404 705458
rect 414804 668454 415404 705222
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 632454 415404 667898
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 596454 415404 631898
rect 414804 596218 414986 596454
rect 415222 596218 415404 596454
rect 414804 596134 415404 596218
rect 414804 595898 414986 596134
rect 415222 595898 415404 596134
rect 414804 584916 415404 595898
rect 432804 704838 433404 705800
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 614454 433404 649898
rect 432804 614218 432986 614454
rect 433222 614218 433404 614454
rect 432804 614134 433404 614218
rect 432804 613898 432986 614134
rect 433222 613898 433404 614134
rect 432804 584916 433404 613898
rect 450804 705778 451404 705800
rect 450804 705542 450986 705778
rect 451222 705542 451404 705778
rect 450804 705458 451404 705542
rect 450804 705222 450986 705458
rect 451222 705222 451404 705458
rect 450804 668454 451404 705222
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 632454 451404 667898
rect 450804 632218 450986 632454
rect 451222 632218 451404 632454
rect 450804 632134 451404 632218
rect 450804 631898 450986 632134
rect 451222 631898 451404 632134
rect 450804 596454 451404 631898
rect 450804 596218 450986 596454
rect 451222 596218 451404 596454
rect 450804 596134 451404 596218
rect 450804 595898 450986 596134
rect 451222 595898 451404 596134
rect 450804 584916 451404 595898
rect 468804 704838 469404 705800
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 650454 469404 685898
rect 468804 650218 468986 650454
rect 469222 650218 469404 650454
rect 468804 650134 469404 650218
rect 468804 649898 468986 650134
rect 469222 649898 469404 650134
rect 468804 614454 469404 649898
rect 468804 614218 468986 614454
rect 469222 614218 469404 614454
rect 468804 614134 469404 614218
rect 468804 613898 468986 614134
rect 469222 613898 469404 614134
rect 468804 584916 469404 613898
rect 486804 705778 487404 705800
rect 486804 705542 486986 705778
rect 487222 705542 487404 705778
rect 486804 705458 487404 705542
rect 486804 705222 486986 705458
rect 487222 705222 487404 705458
rect 486804 668454 487404 705222
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 632454 487404 667898
rect 486804 632218 486986 632454
rect 487222 632218 487404 632454
rect 486804 632134 487404 632218
rect 486804 631898 486986 632134
rect 487222 631898 487404 632134
rect 486804 596454 487404 631898
rect 486804 596218 486986 596454
rect 487222 596218 487404 596454
rect 486804 596134 487404 596218
rect 486804 595898 486986 596134
rect 487222 595898 487404 596134
rect 486804 584916 487404 595898
rect 504804 704838 505404 705800
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 650454 505404 685898
rect 504804 650218 504986 650454
rect 505222 650218 505404 650454
rect 504804 650134 505404 650218
rect 504804 649898 504986 650134
rect 505222 649898 505404 650134
rect 504804 614454 505404 649898
rect 504804 614218 504986 614454
rect 505222 614218 505404 614454
rect 504804 614134 505404 614218
rect 504804 613898 504986 614134
rect 505222 613898 505404 614134
rect 504804 584916 505404 613898
rect 522804 705778 523404 705800
rect 522804 705542 522986 705778
rect 523222 705542 523404 705778
rect 522804 705458 523404 705542
rect 522804 705222 522986 705458
rect 523222 705222 523404 705458
rect 522804 668454 523404 705222
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522804 584916 523404 595898
rect 540804 704838 541404 705800
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 584916 541404 613898
rect 558804 705778 559404 705800
rect 558804 705542 558986 705778
rect 559222 705542 559404 705778
rect 558804 705458 559404 705542
rect 558804 705222 558986 705458
rect 559222 705222 559404 705458
rect 558804 668454 559404 705222
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 584916 559404 595898
rect 576804 704838 577404 705800
rect 586260 705778 586860 705800
rect 586260 705542 586442 705778
rect 586678 705542 586860 705778
rect 586260 705458 586860 705542
rect 586260 705222 586442 705458
rect 586678 705222 586860 705458
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 339216 578454 339536 578476
rect 339216 578218 339258 578454
rect 339494 578218 339536 578454
rect 339216 578134 339536 578218
rect 339216 577898 339258 578134
rect 339494 577898 339536 578134
rect 339216 577876 339536 577898
rect 369936 578454 370256 578476
rect 369936 578218 369978 578454
rect 370214 578218 370256 578454
rect 369936 578134 370256 578218
rect 369936 577898 369978 578134
rect 370214 577898 370256 578134
rect 369936 577876 370256 577898
rect 400656 578454 400976 578476
rect 400656 578218 400698 578454
rect 400934 578218 400976 578454
rect 400656 578134 400976 578218
rect 400656 577898 400698 578134
rect 400934 577898 400976 578134
rect 400656 577876 400976 577898
rect 431376 578454 431696 578476
rect 431376 578218 431418 578454
rect 431654 578218 431696 578454
rect 431376 578134 431696 578218
rect 431376 577898 431418 578134
rect 431654 577898 431696 578134
rect 431376 577876 431696 577898
rect 462096 578454 462416 578476
rect 462096 578218 462138 578454
rect 462374 578218 462416 578454
rect 462096 578134 462416 578218
rect 462096 577898 462138 578134
rect 462374 577898 462416 578134
rect 462096 577876 462416 577898
rect 492816 578454 493136 578476
rect 492816 578218 492858 578454
rect 493094 578218 493136 578454
rect 492816 578134 493136 578218
rect 492816 577898 492858 578134
rect 493094 577898 493136 578134
rect 492816 577876 493136 577898
rect 523536 578454 523856 578476
rect 523536 578218 523578 578454
rect 523814 578218 523856 578454
rect 523536 578134 523856 578218
rect 523536 577898 523578 578134
rect 523814 577898 523856 578134
rect 523536 577876 523856 577898
rect 554256 578454 554576 578476
rect 554256 578218 554298 578454
rect 554534 578218 554576 578454
rect 554256 578134 554576 578218
rect 554256 577898 554298 578134
rect 554534 577898 554576 578134
rect 554256 577876 554576 577898
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 306804 560218 306986 560454
rect 307222 560218 307404 560454
rect 306804 560134 307404 560218
rect 306804 559898 306986 560134
rect 307222 559898 307404 560134
rect 306804 524454 307404 559898
rect 323856 560454 324176 560476
rect 323856 560218 323898 560454
rect 324134 560218 324176 560454
rect 323856 560134 324176 560218
rect 323856 559898 323898 560134
rect 324134 559898 324176 560134
rect 323856 559876 324176 559898
rect 354576 560454 354896 560476
rect 354576 560218 354618 560454
rect 354854 560218 354896 560454
rect 354576 560134 354896 560218
rect 354576 559898 354618 560134
rect 354854 559898 354896 560134
rect 354576 559876 354896 559898
rect 385296 560454 385616 560476
rect 385296 560218 385338 560454
rect 385574 560218 385616 560454
rect 385296 560134 385616 560218
rect 385296 559898 385338 560134
rect 385574 559898 385616 560134
rect 385296 559876 385616 559898
rect 416016 560454 416336 560476
rect 416016 560218 416058 560454
rect 416294 560218 416336 560454
rect 416016 560134 416336 560218
rect 416016 559898 416058 560134
rect 416294 559898 416336 560134
rect 416016 559876 416336 559898
rect 446736 560454 447056 560476
rect 446736 560218 446778 560454
rect 447014 560218 447056 560454
rect 446736 560134 447056 560218
rect 446736 559898 446778 560134
rect 447014 559898 447056 560134
rect 446736 559876 447056 559898
rect 477456 560454 477776 560476
rect 477456 560218 477498 560454
rect 477734 560218 477776 560454
rect 477456 560134 477776 560218
rect 477456 559898 477498 560134
rect 477734 559898 477776 560134
rect 477456 559876 477776 559898
rect 508176 560454 508496 560476
rect 508176 560218 508218 560454
rect 508454 560218 508496 560454
rect 508176 560134 508496 560218
rect 508176 559898 508218 560134
rect 508454 559898 508496 560134
rect 508176 559876 508496 559898
rect 538896 560454 539216 560476
rect 538896 560218 538938 560454
rect 539174 560218 539216 560454
rect 538896 560134 539216 560218
rect 538896 559898 538938 560134
rect 539174 559898 539216 560134
rect 538896 559876 539216 559898
rect 339216 542454 339536 542476
rect 339216 542218 339258 542454
rect 339494 542218 339536 542454
rect 339216 542134 339536 542218
rect 339216 541898 339258 542134
rect 339494 541898 339536 542134
rect 339216 541876 339536 541898
rect 369936 542454 370256 542476
rect 369936 542218 369978 542454
rect 370214 542218 370256 542454
rect 369936 542134 370256 542218
rect 369936 541898 369978 542134
rect 370214 541898 370256 542134
rect 369936 541876 370256 541898
rect 400656 542454 400976 542476
rect 400656 542218 400698 542454
rect 400934 542218 400976 542454
rect 400656 542134 400976 542218
rect 400656 541898 400698 542134
rect 400934 541898 400976 542134
rect 400656 541876 400976 541898
rect 431376 542454 431696 542476
rect 431376 542218 431418 542454
rect 431654 542218 431696 542454
rect 431376 542134 431696 542218
rect 431376 541898 431418 542134
rect 431654 541898 431696 542134
rect 431376 541876 431696 541898
rect 462096 542454 462416 542476
rect 462096 542218 462138 542454
rect 462374 542218 462416 542454
rect 462096 542134 462416 542218
rect 462096 541898 462138 542134
rect 462374 541898 462416 542134
rect 462096 541876 462416 541898
rect 492816 542454 493136 542476
rect 492816 542218 492858 542454
rect 493094 542218 493136 542454
rect 492816 542134 493136 542218
rect 492816 541898 492858 542134
rect 493094 541898 493136 542134
rect 492816 541876 493136 541898
rect 523536 542454 523856 542476
rect 523536 542218 523578 542454
rect 523814 542218 523856 542454
rect 523536 542134 523856 542218
rect 523536 541898 523578 542134
rect 523814 541898 523856 542134
rect 523536 541876 523856 541898
rect 554256 542454 554576 542476
rect 554256 542218 554298 542454
rect 554534 542218 554576 542454
rect 554256 542134 554576 542218
rect 554256 541898 554298 542134
rect 554534 541898 554576 542134
rect 554256 541876 554576 541898
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 306804 524218 306986 524454
rect 307222 524218 307404 524454
rect 306804 524134 307404 524218
rect 306804 523898 306986 524134
rect 307222 523898 307404 524134
rect 306804 488454 307404 523898
rect 323856 524454 324176 524476
rect 323856 524218 323898 524454
rect 324134 524218 324176 524454
rect 323856 524134 324176 524218
rect 323856 523898 323898 524134
rect 324134 523898 324176 524134
rect 323856 523876 324176 523898
rect 354576 524454 354896 524476
rect 354576 524218 354618 524454
rect 354854 524218 354896 524454
rect 354576 524134 354896 524218
rect 354576 523898 354618 524134
rect 354854 523898 354896 524134
rect 354576 523876 354896 523898
rect 385296 524454 385616 524476
rect 385296 524218 385338 524454
rect 385574 524218 385616 524454
rect 385296 524134 385616 524218
rect 385296 523898 385338 524134
rect 385574 523898 385616 524134
rect 385296 523876 385616 523898
rect 416016 524454 416336 524476
rect 416016 524218 416058 524454
rect 416294 524218 416336 524454
rect 416016 524134 416336 524218
rect 416016 523898 416058 524134
rect 416294 523898 416336 524134
rect 416016 523876 416336 523898
rect 446736 524454 447056 524476
rect 446736 524218 446778 524454
rect 447014 524218 447056 524454
rect 446736 524134 447056 524218
rect 446736 523898 446778 524134
rect 447014 523898 447056 524134
rect 446736 523876 447056 523898
rect 477456 524454 477776 524476
rect 477456 524218 477498 524454
rect 477734 524218 477776 524454
rect 477456 524134 477776 524218
rect 477456 523898 477498 524134
rect 477734 523898 477776 524134
rect 477456 523876 477776 523898
rect 508176 524454 508496 524476
rect 508176 524218 508218 524454
rect 508454 524218 508496 524454
rect 508176 524134 508496 524218
rect 508176 523898 508218 524134
rect 508454 523898 508496 524134
rect 508176 523876 508496 523898
rect 538896 524454 539216 524476
rect 538896 524218 538938 524454
rect 539174 524218 539216 524454
rect 538896 524134 539216 524218
rect 538896 523898 538938 524134
rect 539174 523898 539216 524134
rect 538896 523876 539216 523898
rect 339216 506454 339536 506476
rect 339216 506218 339258 506454
rect 339494 506218 339536 506454
rect 339216 506134 339536 506218
rect 339216 505898 339258 506134
rect 339494 505898 339536 506134
rect 339216 505876 339536 505898
rect 369936 506454 370256 506476
rect 369936 506218 369978 506454
rect 370214 506218 370256 506454
rect 369936 506134 370256 506218
rect 369936 505898 369978 506134
rect 370214 505898 370256 506134
rect 369936 505876 370256 505898
rect 400656 506454 400976 506476
rect 400656 506218 400698 506454
rect 400934 506218 400976 506454
rect 400656 506134 400976 506218
rect 400656 505898 400698 506134
rect 400934 505898 400976 506134
rect 400656 505876 400976 505898
rect 431376 506454 431696 506476
rect 431376 506218 431418 506454
rect 431654 506218 431696 506454
rect 431376 506134 431696 506218
rect 431376 505898 431418 506134
rect 431654 505898 431696 506134
rect 431376 505876 431696 505898
rect 462096 506454 462416 506476
rect 462096 506218 462138 506454
rect 462374 506218 462416 506454
rect 462096 506134 462416 506218
rect 462096 505898 462138 506134
rect 462374 505898 462416 506134
rect 462096 505876 462416 505898
rect 492816 506454 493136 506476
rect 492816 506218 492858 506454
rect 493094 506218 493136 506454
rect 492816 506134 493136 506218
rect 492816 505898 492858 506134
rect 493094 505898 493136 506134
rect 492816 505876 493136 505898
rect 523536 506454 523856 506476
rect 523536 506218 523578 506454
rect 523814 506218 523856 506454
rect 523536 506134 523856 506218
rect 523536 505898 523578 506134
rect 523814 505898 523856 506134
rect 523536 505876 523856 505898
rect 554256 506454 554576 506476
rect 554256 506218 554298 506454
rect 554534 506218 554576 506454
rect 554256 506134 554576 506218
rect 554256 505898 554298 506134
rect 554534 505898 554576 506134
rect 554256 505876 554576 505898
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 306804 488218 306986 488454
rect 307222 488218 307404 488454
rect 306804 488134 307404 488218
rect 306804 487898 306986 488134
rect 307222 487898 307404 488134
rect 306804 452454 307404 487898
rect 323856 488454 324176 488476
rect 323856 488218 323898 488454
rect 324134 488218 324176 488454
rect 323856 488134 324176 488218
rect 323856 487898 323898 488134
rect 324134 487898 324176 488134
rect 323856 487876 324176 487898
rect 354576 488454 354896 488476
rect 354576 488218 354618 488454
rect 354854 488218 354896 488454
rect 354576 488134 354896 488218
rect 354576 487898 354618 488134
rect 354854 487898 354896 488134
rect 354576 487876 354896 487898
rect 385296 488454 385616 488476
rect 385296 488218 385338 488454
rect 385574 488218 385616 488454
rect 385296 488134 385616 488218
rect 385296 487898 385338 488134
rect 385574 487898 385616 488134
rect 385296 487876 385616 487898
rect 416016 488454 416336 488476
rect 416016 488218 416058 488454
rect 416294 488218 416336 488454
rect 416016 488134 416336 488218
rect 416016 487898 416058 488134
rect 416294 487898 416336 488134
rect 416016 487876 416336 487898
rect 446736 488454 447056 488476
rect 446736 488218 446778 488454
rect 447014 488218 447056 488454
rect 446736 488134 447056 488218
rect 446736 487898 446778 488134
rect 447014 487898 447056 488134
rect 446736 487876 447056 487898
rect 477456 488454 477776 488476
rect 477456 488218 477498 488454
rect 477734 488218 477776 488454
rect 477456 488134 477776 488218
rect 477456 487898 477498 488134
rect 477734 487898 477776 488134
rect 477456 487876 477776 487898
rect 508176 488454 508496 488476
rect 508176 488218 508218 488454
rect 508454 488218 508496 488454
rect 508176 488134 508496 488218
rect 508176 487898 508218 488134
rect 508454 487898 508496 488134
rect 508176 487876 508496 487898
rect 538896 488454 539216 488476
rect 538896 488218 538938 488454
rect 539174 488218 539216 488454
rect 538896 488134 539216 488218
rect 538896 487898 538938 488134
rect 539174 487898 539216 488134
rect 538896 487876 539216 487898
rect 339216 470454 339536 470476
rect 339216 470218 339258 470454
rect 339494 470218 339536 470454
rect 339216 470134 339536 470218
rect 339216 469898 339258 470134
rect 339494 469898 339536 470134
rect 339216 469876 339536 469898
rect 369936 470454 370256 470476
rect 369936 470218 369978 470454
rect 370214 470218 370256 470454
rect 369936 470134 370256 470218
rect 369936 469898 369978 470134
rect 370214 469898 370256 470134
rect 369936 469876 370256 469898
rect 400656 470454 400976 470476
rect 400656 470218 400698 470454
rect 400934 470218 400976 470454
rect 400656 470134 400976 470218
rect 400656 469898 400698 470134
rect 400934 469898 400976 470134
rect 400656 469876 400976 469898
rect 431376 470454 431696 470476
rect 431376 470218 431418 470454
rect 431654 470218 431696 470454
rect 431376 470134 431696 470218
rect 431376 469898 431418 470134
rect 431654 469898 431696 470134
rect 431376 469876 431696 469898
rect 462096 470454 462416 470476
rect 462096 470218 462138 470454
rect 462374 470218 462416 470454
rect 462096 470134 462416 470218
rect 462096 469898 462138 470134
rect 462374 469898 462416 470134
rect 462096 469876 462416 469898
rect 492816 470454 493136 470476
rect 492816 470218 492858 470454
rect 493094 470218 493136 470454
rect 492816 470134 493136 470218
rect 492816 469898 492858 470134
rect 493094 469898 493136 470134
rect 492816 469876 493136 469898
rect 523536 470454 523856 470476
rect 523536 470218 523578 470454
rect 523814 470218 523856 470454
rect 523536 470134 523856 470218
rect 523536 469898 523578 470134
rect 523814 469898 523856 470134
rect 523536 469876 523856 469898
rect 554256 470454 554576 470476
rect 554256 470218 554298 470454
rect 554534 470218 554576 470454
rect 554256 470134 554576 470218
rect 554256 469898 554298 470134
rect 554534 469898 554576 470134
rect 554256 469876 554576 469898
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 306804 452218 306986 452454
rect 307222 452218 307404 452454
rect 306804 452134 307404 452218
rect 306804 451898 306986 452134
rect 307222 451898 307404 452134
rect 306804 416454 307404 451898
rect 323856 452454 324176 452476
rect 323856 452218 323898 452454
rect 324134 452218 324176 452454
rect 323856 452134 324176 452218
rect 323856 451898 323898 452134
rect 324134 451898 324176 452134
rect 323856 451876 324176 451898
rect 354576 452454 354896 452476
rect 354576 452218 354618 452454
rect 354854 452218 354896 452454
rect 354576 452134 354896 452218
rect 354576 451898 354618 452134
rect 354854 451898 354896 452134
rect 354576 451876 354896 451898
rect 385296 452454 385616 452476
rect 385296 452218 385338 452454
rect 385574 452218 385616 452454
rect 385296 452134 385616 452218
rect 385296 451898 385338 452134
rect 385574 451898 385616 452134
rect 385296 451876 385616 451898
rect 416016 452454 416336 452476
rect 416016 452218 416058 452454
rect 416294 452218 416336 452454
rect 416016 452134 416336 452218
rect 416016 451898 416058 452134
rect 416294 451898 416336 452134
rect 416016 451876 416336 451898
rect 446736 452454 447056 452476
rect 446736 452218 446778 452454
rect 447014 452218 447056 452454
rect 446736 452134 447056 452218
rect 446736 451898 446778 452134
rect 447014 451898 447056 452134
rect 446736 451876 447056 451898
rect 477456 452454 477776 452476
rect 477456 452218 477498 452454
rect 477734 452218 477776 452454
rect 477456 452134 477776 452218
rect 477456 451898 477498 452134
rect 477734 451898 477776 452134
rect 477456 451876 477776 451898
rect 508176 452454 508496 452476
rect 508176 452218 508218 452454
rect 508454 452218 508496 452454
rect 508176 452134 508496 452218
rect 508176 451898 508218 452134
rect 508454 451898 508496 452134
rect 508176 451876 508496 451898
rect 538896 452454 539216 452476
rect 538896 452218 538938 452454
rect 539174 452218 539216 452454
rect 538896 452134 539216 452218
rect 538896 451898 538938 452134
rect 539174 451898 539216 452134
rect 538896 451876 539216 451898
rect 339216 434454 339536 434476
rect 339216 434218 339258 434454
rect 339494 434218 339536 434454
rect 339216 434134 339536 434218
rect 339216 433898 339258 434134
rect 339494 433898 339536 434134
rect 339216 433876 339536 433898
rect 369936 434454 370256 434476
rect 369936 434218 369978 434454
rect 370214 434218 370256 434454
rect 369936 434134 370256 434218
rect 369936 433898 369978 434134
rect 370214 433898 370256 434134
rect 369936 433876 370256 433898
rect 400656 434454 400976 434476
rect 400656 434218 400698 434454
rect 400934 434218 400976 434454
rect 400656 434134 400976 434218
rect 400656 433898 400698 434134
rect 400934 433898 400976 434134
rect 400656 433876 400976 433898
rect 431376 434454 431696 434476
rect 431376 434218 431418 434454
rect 431654 434218 431696 434454
rect 431376 434134 431696 434218
rect 431376 433898 431418 434134
rect 431654 433898 431696 434134
rect 431376 433876 431696 433898
rect 462096 434454 462416 434476
rect 462096 434218 462138 434454
rect 462374 434218 462416 434454
rect 462096 434134 462416 434218
rect 462096 433898 462138 434134
rect 462374 433898 462416 434134
rect 462096 433876 462416 433898
rect 492816 434454 493136 434476
rect 492816 434218 492858 434454
rect 493094 434218 493136 434454
rect 492816 434134 493136 434218
rect 492816 433898 492858 434134
rect 493094 433898 493136 434134
rect 492816 433876 493136 433898
rect 523536 434454 523856 434476
rect 523536 434218 523578 434454
rect 523814 434218 523856 434454
rect 523536 434134 523856 434218
rect 523536 433898 523578 434134
rect 523814 433898 523856 434134
rect 523536 433876 523856 433898
rect 554256 434454 554576 434476
rect 554256 434218 554298 434454
rect 554534 434218 554576 434454
rect 554256 434134 554576 434218
rect 554256 433898 554298 434134
rect 554534 433898 554576 434134
rect 554256 433876 554576 433898
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 306804 416218 306986 416454
rect 307222 416218 307404 416454
rect 306804 416134 307404 416218
rect 306804 415898 306986 416134
rect 307222 415898 307404 416134
rect 306804 380454 307404 415898
rect 323856 416454 324176 416476
rect 323856 416218 323898 416454
rect 324134 416218 324176 416454
rect 323856 416134 324176 416218
rect 323856 415898 323898 416134
rect 324134 415898 324176 416134
rect 323856 415876 324176 415898
rect 354576 416454 354896 416476
rect 354576 416218 354618 416454
rect 354854 416218 354896 416454
rect 354576 416134 354896 416218
rect 354576 415898 354618 416134
rect 354854 415898 354896 416134
rect 354576 415876 354896 415898
rect 385296 416454 385616 416476
rect 385296 416218 385338 416454
rect 385574 416218 385616 416454
rect 385296 416134 385616 416218
rect 385296 415898 385338 416134
rect 385574 415898 385616 416134
rect 385296 415876 385616 415898
rect 416016 416454 416336 416476
rect 416016 416218 416058 416454
rect 416294 416218 416336 416454
rect 416016 416134 416336 416218
rect 416016 415898 416058 416134
rect 416294 415898 416336 416134
rect 416016 415876 416336 415898
rect 446736 416454 447056 416476
rect 446736 416218 446778 416454
rect 447014 416218 447056 416454
rect 446736 416134 447056 416218
rect 446736 415898 446778 416134
rect 447014 415898 447056 416134
rect 446736 415876 447056 415898
rect 477456 416454 477776 416476
rect 477456 416218 477498 416454
rect 477734 416218 477776 416454
rect 477456 416134 477776 416218
rect 477456 415898 477498 416134
rect 477734 415898 477776 416134
rect 477456 415876 477776 415898
rect 508176 416454 508496 416476
rect 508176 416218 508218 416454
rect 508454 416218 508496 416454
rect 508176 416134 508496 416218
rect 508176 415898 508218 416134
rect 508454 415898 508496 416134
rect 508176 415876 508496 415898
rect 538896 416454 539216 416476
rect 538896 416218 538938 416454
rect 539174 416218 539216 416454
rect 538896 416134 539216 416218
rect 538896 415898 538938 416134
rect 539174 415898 539216 416134
rect 538896 415876 539216 415898
rect 339216 398454 339536 398476
rect 339216 398218 339258 398454
rect 339494 398218 339536 398454
rect 339216 398134 339536 398218
rect 339216 397898 339258 398134
rect 339494 397898 339536 398134
rect 339216 397876 339536 397898
rect 369936 398454 370256 398476
rect 369936 398218 369978 398454
rect 370214 398218 370256 398454
rect 369936 398134 370256 398218
rect 369936 397898 369978 398134
rect 370214 397898 370256 398134
rect 369936 397876 370256 397898
rect 400656 398454 400976 398476
rect 400656 398218 400698 398454
rect 400934 398218 400976 398454
rect 400656 398134 400976 398218
rect 400656 397898 400698 398134
rect 400934 397898 400976 398134
rect 400656 397876 400976 397898
rect 431376 398454 431696 398476
rect 431376 398218 431418 398454
rect 431654 398218 431696 398454
rect 431376 398134 431696 398218
rect 431376 397898 431418 398134
rect 431654 397898 431696 398134
rect 431376 397876 431696 397898
rect 462096 398454 462416 398476
rect 462096 398218 462138 398454
rect 462374 398218 462416 398454
rect 462096 398134 462416 398218
rect 462096 397898 462138 398134
rect 462374 397898 462416 398134
rect 462096 397876 462416 397898
rect 492816 398454 493136 398476
rect 492816 398218 492858 398454
rect 493094 398218 493136 398454
rect 492816 398134 493136 398218
rect 492816 397898 492858 398134
rect 493094 397898 493136 398134
rect 492816 397876 493136 397898
rect 523536 398454 523856 398476
rect 523536 398218 523578 398454
rect 523814 398218 523856 398454
rect 523536 398134 523856 398218
rect 523536 397898 523578 398134
rect 523814 397898 523856 398134
rect 523536 397876 523856 397898
rect 554256 398454 554576 398476
rect 554256 398218 554298 398454
rect 554534 398218 554576 398454
rect 554256 398134 554576 398218
rect 554256 397898 554298 398134
rect 554534 397898 554576 398134
rect 554256 397876 554576 397898
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 306804 380218 306986 380454
rect 307222 380218 307404 380454
rect 306804 380134 307404 380218
rect 306804 379898 306986 380134
rect 307222 379898 307404 380134
rect 306804 356560 307404 379898
rect 324804 362454 325404 382916
rect 324804 362218 324986 362454
rect 325222 362218 325404 362454
rect 324804 362134 325404 362218
rect 324804 361898 324986 362134
rect 325222 361898 325404 362134
rect 292112 344454 292432 344476
rect 292112 344218 292154 344454
rect 292390 344218 292432 344454
rect 292112 344134 292432 344218
rect 292112 343898 292154 344134
rect 292390 343898 292432 344134
rect 292112 343876 292432 343898
rect 252804 326218 252986 326454
rect 253222 326218 253404 326454
rect 252804 326134 253404 326218
rect 252804 325898 252986 326134
rect 253222 325898 253404 326134
rect 252804 290454 253404 325898
rect 276752 326454 277072 326476
rect 276752 326218 276794 326454
rect 277030 326218 277072 326454
rect 276752 326134 277072 326218
rect 276752 325898 276794 326134
rect 277030 325898 277072 326134
rect 276752 325876 277072 325898
rect 307472 326454 307792 326476
rect 307472 326218 307514 326454
rect 307750 326218 307792 326454
rect 307472 326134 307792 326218
rect 307472 325898 307514 326134
rect 307750 325898 307792 326134
rect 307472 325876 307792 325898
rect 324804 326454 325404 361898
rect 324804 326218 324986 326454
rect 325222 326218 325404 326454
rect 324804 326134 325404 326218
rect 324804 325898 324986 326134
rect 325222 325898 325404 326134
rect 252804 290218 252986 290454
rect 253222 290218 253404 290454
rect 252804 290134 253404 290218
rect 252804 289898 252986 290134
rect 253222 289898 253404 290134
rect 252804 274600 253404 289898
rect 270804 308454 271404 314560
rect 270804 308218 270986 308454
rect 271222 308218 271404 308454
rect 270804 308134 271404 308218
rect 270804 307898 270986 308134
rect 271222 307898 271404 308134
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 270804 272454 271404 307898
rect 270804 272218 270986 272454
rect 271222 272218 271404 272454
rect 270804 272134 271404 272218
rect 270804 271898 270986 272134
rect 271222 271898 271404 272134
rect 47088 254454 47408 254476
rect 47088 254218 47130 254454
rect 47366 254218 47408 254454
rect 47088 254134 47408 254218
rect 47088 253898 47130 254134
rect 47366 253898 47408 254134
rect 47088 253876 47408 253898
rect 77808 254454 78128 254476
rect 77808 254218 77850 254454
rect 78086 254218 78128 254454
rect 77808 254134 78128 254218
rect 77808 253898 77850 254134
rect 78086 253898 78128 254134
rect 77808 253876 78128 253898
rect 108528 254454 108848 254476
rect 108528 254218 108570 254454
rect 108806 254218 108848 254454
rect 108528 254134 108848 254218
rect 108528 253898 108570 254134
rect 108806 253898 108848 254134
rect 108528 253876 108848 253898
rect 139248 254454 139568 254476
rect 139248 254218 139290 254454
rect 139526 254218 139568 254454
rect 139248 254134 139568 254218
rect 139248 253898 139290 254134
rect 139526 253898 139568 254134
rect 139248 253876 139568 253898
rect 169968 254454 170288 254476
rect 169968 254218 170010 254454
rect 170246 254218 170288 254454
rect 169968 254134 170288 254218
rect 169968 253898 170010 254134
rect 170246 253898 170288 254134
rect 169968 253876 170288 253898
rect 200688 254454 201008 254476
rect 200688 254218 200730 254454
rect 200966 254218 201008 254454
rect 200688 254134 201008 254218
rect 200688 253898 200730 254134
rect 200966 253898 201008 254134
rect 200688 253876 201008 253898
rect 231408 254454 231728 254476
rect 231408 254218 231450 254454
rect 231686 254218 231728 254454
rect 231408 254134 231728 254218
rect 231408 253898 231450 254134
rect 231686 253898 231728 254134
rect 231408 253876 231728 253898
rect 262128 254454 262448 254476
rect 262128 254218 262170 254454
rect 262406 254218 262448 254454
rect 262128 254134 262448 254218
rect 262128 253898 262170 254134
rect 262406 253898 262448 254134
rect 262128 253876 262448 253898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 31728 236454 32048 236476
rect 31728 236218 31770 236454
rect 32006 236218 32048 236454
rect 31728 236134 32048 236218
rect 31728 235898 31770 236134
rect 32006 235898 32048 236134
rect 31728 235876 32048 235898
rect 62448 236454 62768 236476
rect 62448 236218 62490 236454
rect 62726 236218 62768 236454
rect 62448 236134 62768 236218
rect 62448 235898 62490 236134
rect 62726 235898 62768 236134
rect 62448 235876 62768 235898
rect 93168 236454 93488 236476
rect 93168 236218 93210 236454
rect 93446 236218 93488 236454
rect 93168 236134 93488 236218
rect 93168 235898 93210 236134
rect 93446 235898 93488 236134
rect 93168 235876 93488 235898
rect 123888 236454 124208 236476
rect 123888 236218 123930 236454
rect 124166 236218 124208 236454
rect 123888 236134 124208 236218
rect 123888 235898 123930 236134
rect 124166 235898 124208 236134
rect 123888 235876 124208 235898
rect 154608 236454 154928 236476
rect 154608 236218 154650 236454
rect 154886 236218 154928 236454
rect 154608 236134 154928 236218
rect 154608 235898 154650 236134
rect 154886 235898 154928 236134
rect 154608 235876 154928 235898
rect 185328 236454 185648 236476
rect 185328 236218 185370 236454
rect 185606 236218 185648 236454
rect 185328 236134 185648 236218
rect 185328 235898 185370 236134
rect 185606 235898 185648 236134
rect 185328 235876 185648 235898
rect 216048 236454 216368 236476
rect 216048 236218 216090 236454
rect 216326 236218 216368 236454
rect 216048 236134 216368 236218
rect 216048 235898 216090 236134
rect 216326 235898 216368 236134
rect 216048 235876 216368 235898
rect 246768 236454 247088 236476
rect 246768 236218 246810 236454
rect 247046 236218 247088 236454
rect 246768 236134 247088 236218
rect 246768 235898 246810 236134
rect 247046 235898 247088 236134
rect 246768 235876 247088 235898
rect 270804 236454 271404 271898
rect 270804 236218 270986 236454
rect 271222 236218 271404 236454
rect 270804 236134 271404 236218
rect 270804 235898 270986 236134
rect 271222 235898 271404 236134
rect 47088 218454 47408 218476
rect 47088 218218 47130 218454
rect 47366 218218 47408 218454
rect 47088 218134 47408 218218
rect 47088 217898 47130 218134
rect 47366 217898 47408 218134
rect 47088 217876 47408 217898
rect 77808 218454 78128 218476
rect 77808 218218 77850 218454
rect 78086 218218 78128 218454
rect 77808 218134 78128 218218
rect 77808 217898 77850 218134
rect 78086 217898 78128 218134
rect 77808 217876 78128 217898
rect 108528 218454 108848 218476
rect 108528 218218 108570 218454
rect 108806 218218 108848 218454
rect 108528 218134 108848 218218
rect 108528 217898 108570 218134
rect 108806 217898 108848 218134
rect 108528 217876 108848 217898
rect 139248 218454 139568 218476
rect 139248 218218 139290 218454
rect 139526 218218 139568 218454
rect 139248 218134 139568 218218
rect 139248 217898 139290 218134
rect 139526 217898 139568 218134
rect 139248 217876 139568 217898
rect 169968 218454 170288 218476
rect 169968 218218 170010 218454
rect 170246 218218 170288 218454
rect 169968 218134 170288 218218
rect 169968 217898 170010 218134
rect 170246 217898 170288 218134
rect 169968 217876 170288 217898
rect 200688 218454 201008 218476
rect 200688 218218 200730 218454
rect 200966 218218 201008 218454
rect 200688 218134 201008 218218
rect 200688 217898 200730 218134
rect 200966 217898 201008 218134
rect 200688 217876 201008 217898
rect 231408 218454 231728 218476
rect 231408 218218 231450 218454
rect 231686 218218 231728 218454
rect 231408 218134 231728 218218
rect 231408 217898 231450 218134
rect 231686 217898 231728 218134
rect 231408 217876 231728 217898
rect 262128 218454 262448 218476
rect 262128 218218 262170 218454
rect 262406 218218 262448 218454
rect 262128 218134 262448 218218
rect 262128 217898 262170 218134
rect 262406 217898 262448 218134
rect 262128 217876 262448 217898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 31728 200454 32048 200476
rect 31728 200218 31770 200454
rect 32006 200218 32048 200454
rect 31728 200134 32048 200218
rect 31728 199898 31770 200134
rect 32006 199898 32048 200134
rect 31728 199876 32048 199898
rect 62448 200454 62768 200476
rect 62448 200218 62490 200454
rect 62726 200218 62768 200454
rect 62448 200134 62768 200218
rect 62448 199898 62490 200134
rect 62726 199898 62768 200134
rect 62448 199876 62768 199898
rect 93168 200454 93488 200476
rect 93168 200218 93210 200454
rect 93446 200218 93488 200454
rect 93168 200134 93488 200218
rect 93168 199898 93210 200134
rect 93446 199898 93488 200134
rect 93168 199876 93488 199898
rect 123888 200454 124208 200476
rect 123888 200218 123930 200454
rect 124166 200218 124208 200454
rect 123888 200134 124208 200218
rect 123888 199898 123930 200134
rect 124166 199898 124208 200134
rect 123888 199876 124208 199898
rect 154608 200454 154928 200476
rect 154608 200218 154650 200454
rect 154886 200218 154928 200454
rect 154608 200134 154928 200218
rect 154608 199898 154650 200134
rect 154886 199898 154928 200134
rect 154608 199876 154928 199898
rect 185328 200454 185648 200476
rect 185328 200218 185370 200454
rect 185606 200218 185648 200454
rect 185328 200134 185648 200218
rect 185328 199898 185370 200134
rect 185606 199898 185648 200134
rect 185328 199876 185648 199898
rect 216048 200454 216368 200476
rect 216048 200218 216090 200454
rect 216326 200218 216368 200454
rect 216048 200134 216368 200218
rect 216048 199898 216090 200134
rect 216326 199898 216368 200134
rect 216048 199876 216368 199898
rect 246768 200454 247088 200476
rect 246768 200218 246810 200454
rect 247046 200218 247088 200454
rect 246768 200134 247088 200218
rect 246768 199898 246810 200134
rect 247046 199898 247088 200134
rect 246768 199876 247088 199898
rect 270804 200454 271404 235898
rect 270804 200218 270986 200454
rect 271222 200218 271404 200454
rect 270804 200134 271404 200218
rect 270804 199898 270986 200134
rect 271222 199898 271404 200134
rect 47088 182454 47408 182476
rect 47088 182218 47130 182454
rect 47366 182218 47408 182454
rect 47088 182134 47408 182218
rect 47088 181898 47130 182134
rect 47366 181898 47408 182134
rect 47088 181876 47408 181898
rect 77808 182454 78128 182476
rect 77808 182218 77850 182454
rect 78086 182218 78128 182454
rect 77808 182134 78128 182218
rect 77808 181898 77850 182134
rect 78086 181898 78128 182134
rect 77808 181876 78128 181898
rect 108528 182454 108848 182476
rect 108528 182218 108570 182454
rect 108806 182218 108848 182454
rect 108528 182134 108848 182218
rect 108528 181898 108570 182134
rect 108806 181898 108848 182134
rect 108528 181876 108848 181898
rect 139248 182454 139568 182476
rect 139248 182218 139290 182454
rect 139526 182218 139568 182454
rect 139248 182134 139568 182218
rect 139248 181898 139290 182134
rect 139526 181898 139568 182134
rect 139248 181876 139568 181898
rect 169968 182454 170288 182476
rect 169968 182218 170010 182454
rect 170246 182218 170288 182454
rect 169968 182134 170288 182218
rect 169968 181898 170010 182134
rect 170246 181898 170288 182134
rect 169968 181876 170288 181898
rect 200688 182454 201008 182476
rect 200688 182218 200730 182454
rect 200966 182218 201008 182454
rect 200688 182134 201008 182218
rect 200688 181898 200730 182134
rect 200966 181898 201008 182134
rect 200688 181876 201008 181898
rect 231408 182454 231728 182476
rect 231408 182218 231450 182454
rect 231686 182218 231728 182454
rect 231408 182134 231728 182218
rect 231408 181898 231450 182134
rect 231686 181898 231728 182134
rect 231408 181876 231728 181898
rect 262128 182454 262448 182476
rect 262128 182218 262170 182454
rect 262406 182218 262448 182454
rect 262128 182134 262448 182218
rect 262128 181898 262170 182134
rect 262406 181898 262448 182134
rect 262128 181876 262448 181898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 31728 164454 32048 164476
rect 31728 164218 31770 164454
rect 32006 164218 32048 164454
rect 31728 164134 32048 164218
rect 31728 163898 31770 164134
rect 32006 163898 32048 164134
rect 31728 163876 32048 163898
rect 62448 164454 62768 164476
rect 62448 164218 62490 164454
rect 62726 164218 62768 164454
rect 62448 164134 62768 164218
rect 62448 163898 62490 164134
rect 62726 163898 62768 164134
rect 62448 163876 62768 163898
rect 93168 164454 93488 164476
rect 93168 164218 93210 164454
rect 93446 164218 93488 164454
rect 93168 164134 93488 164218
rect 93168 163898 93210 164134
rect 93446 163898 93488 164134
rect 93168 163876 93488 163898
rect 123888 164454 124208 164476
rect 123888 164218 123930 164454
rect 124166 164218 124208 164454
rect 123888 164134 124208 164218
rect 123888 163898 123930 164134
rect 124166 163898 124208 164134
rect 123888 163876 124208 163898
rect 154608 164454 154928 164476
rect 154608 164218 154650 164454
rect 154886 164218 154928 164454
rect 154608 164134 154928 164218
rect 154608 163898 154650 164134
rect 154886 163898 154928 164134
rect 154608 163876 154928 163898
rect 185328 164454 185648 164476
rect 185328 164218 185370 164454
rect 185606 164218 185648 164454
rect 185328 164134 185648 164218
rect 185328 163898 185370 164134
rect 185606 163898 185648 164134
rect 185328 163876 185648 163898
rect 216048 164454 216368 164476
rect 216048 164218 216090 164454
rect 216326 164218 216368 164454
rect 216048 164134 216368 164218
rect 216048 163898 216090 164134
rect 216326 163898 216368 164134
rect 216048 163876 216368 163898
rect 246768 164454 247088 164476
rect 246768 164218 246810 164454
rect 247046 164218 247088 164454
rect 246768 164134 247088 164218
rect 246768 163898 246810 164134
rect 247046 163898 247088 164134
rect 246768 163876 247088 163898
rect 270804 164454 271404 199898
rect 270804 164218 270986 164454
rect 271222 164218 271404 164454
rect 270804 164134 271404 164218
rect 270804 163898 270986 164134
rect 271222 163898 271404 164134
rect 47088 146454 47408 146476
rect 47088 146218 47130 146454
rect 47366 146218 47408 146454
rect 47088 146134 47408 146218
rect 47088 145898 47130 146134
rect 47366 145898 47408 146134
rect 47088 145876 47408 145898
rect 77808 146454 78128 146476
rect 77808 146218 77850 146454
rect 78086 146218 78128 146454
rect 77808 146134 78128 146218
rect 77808 145898 77850 146134
rect 78086 145898 78128 146134
rect 77808 145876 78128 145898
rect 108528 146454 108848 146476
rect 108528 146218 108570 146454
rect 108806 146218 108848 146454
rect 108528 146134 108848 146218
rect 108528 145898 108570 146134
rect 108806 145898 108848 146134
rect 108528 145876 108848 145898
rect 139248 146454 139568 146476
rect 139248 146218 139290 146454
rect 139526 146218 139568 146454
rect 139248 146134 139568 146218
rect 139248 145898 139290 146134
rect 139526 145898 139568 146134
rect 139248 145876 139568 145898
rect 169968 146454 170288 146476
rect 169968 146218 170010 146454
rect 170246 146218 170288 146454
rect 169968 146134 170288 146218
rect 169968 145898 170010 146134
rect 170246 145898 170288 146134
rect 169968 145876 170288 145898
rect 200688 146454 201008 146476
rect 200688 146218 200730 146454
rect 200966 146218 201008 146454
rect 200688 146134 201008 146218
rect 200688 145898 200730 146134
rect 200966 145898 201008 146134
rect 200688 145876 201008 145898
rect 231408 146454 231728 146476
rect 231408 146218 231450 146454
rect 231686 146218 231728 146454
rect 231408 146134 231728 146218
rect 231408 145898 231450 146134
rect 231686 145898 231728 146134
rect 231408 145876 231728 145898
rect 262128 146454 262448 146476
rect 262128 146218 262170 146454
rect 262406 146218 262448 146454
rect 262128 146134 262448 146218
rect 262128 145898 262170 146134
rect 262406 145898 262448 146134
rect 262128 145876 262448 145898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 31728 128454 32048 128476
rect 31728 128218 31770 128454
rect 32006 128218 32048 128454
rect 31728 128134 32048 128218
rect 31728 127898 31770 128134
rect 32006 127898 32048 128134
rect 31728 127876 32048 127898
rect 62448 128454 62768 128476
rect 62448 128218 62490 128454
rect 62726 128218 62768 128454
rect 62448 128134 62768 128218
rect 62448 127898 62490 128134
rect 62726 127898 62768 128134
rect 62448 127876 62768 127898
rect 93168 128454 93488 128476
rect 93168 128218 93210 128454
rect 93446 128218 93488 128454
rect 93168 128134 93488 128218
rect 93168 127898 93210 128134
rect 93446 127898 93488 128134
rect 93168 127876 93488 127898
rect 123888 128454 124208 128476
rect 123888 128218 123930 128454
rect 124166 128218 124208 128454
rect 123888 128134 124208 128218
rect 123888 127898 123930 128134
rect 124166 127898 124208 128134
rect 123888 127876 124208 127898
rect 154608 128454 154928 128476
rect 154608 128218 154650 128454
rect 154886 128218 154928 128454
rect 154608 128134 154928 128218
rect 154608 127898 154650 128134
rect 154886 127898 154928 128134
rect 154608 127876 154928 127898
rect 185328 128454 185648 128476
rect 185328 128218 185370 128454
rect 185606 128218 185648 128454
rect 185328 128134 185648 128218
rect 185328 127898 185370 128134
rect 185606 127898 185648 128134
rect 185328 127876 185648 127898
rect 216048 128454 216368 128476
rect 216048 128218 216090 128454
rect 216326 128218 216368 128454
rect 216048 128134 216368 128218
rect 216048 127898 216090 128134
rect 216326 127898 216368 128134
rect 216048 127876 216368 127898
rect 246768 128454 247088 128476
rect 246768 128218 246810 128454
rect 247046 128218 247088 128454
rect 246768 128134 247088 128218
rect 246768 127898 246810 128134
rect 247046 127898 247088 128134
rect 246768 127876 247088 127898
rect 270804 128454 271404 163898
rect 270804 128218 270986 128454
rect 271222 128218 271404 128454
rect 270804 128134 271404 128218
rect 270804 127898 270986 128134
rect 271222 127898 271404 128134
rect 47088 110454 47408 110476
rect 47088 110218 47130 110454
rect 47366 110218 47408 110454
rect 47088 110134 47408 110218
rect 47088 109898 47130 110134
rect 47366 109898 47408 110134
rect 47088 109876 47408 109898
rect 77808 110454 78128 110476
rect 77808 110218 77850 110454
rect 78086 110218 78128 110454
rect 77808 110134 78128 110218
rect 77808 109898 77850 110134
rect 78086 109898 78128 110134
rect 77808 109876 78128 109898
rect 108528 110454 108848 110476
rect 108528 110218 108570 110454
rect 108806 110218 108848 110454
rect 108528 110134 108848 110218
rect 108528 109898 108570 110134
rect 108806 109898 108848 110134
rect 108528 109876 108848 109898
rect 139248 110454 139568 110476
rect 139248 110218 139290 110454
rect 139526 110218 139568 110454
rect 139248 110134 139568 110218
rect 139248 109898 139290 110134
rect 139526 109898 139568 110134
rect 139248 109876 139568 109898
rect 169968 110454 170288 110476
rect 169968 110218 170010 110454
rect 170246 110218 170288 110454
rect 169968 110134 170288 110218
rect 169968 109898 170010 110134
rect 170246 109898 170288 110134
rect 169968 109876 170288 109898
rect 200688 110454 201008 110476
rect 200688 110218 200730 110454
rect 200966 110218 201008 110454
rect 200688 110134 201008 110218
rect 200688 109898 200730 110134
rect 200966 109898 201008 110134
rect 200688 109876 201008 109898
rect 231408 110454 231728 110476
rect 231408 110218 231450 110454
rect 231686 110218 231728 110454
rect 231408 110134 231728 110218
rect 231408 109898 231450 110134
rect 231686 109898 231728 110134
rect 231408 109876 231728 109898
rect 262128 110454 262448 110476
rect 262128 110218 262170 110454
rect 262406 110218 262448 110454
rect 262128 110134 262448 110218
rect 262128 109898 262170 110134
rect 262406 109898 262448 110134
rect 262128 109876 262448 109898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 31728 92454 32048 92476
rect 31728 92218 31770 92454
rect 32006 92218 32048 92454
rect 31728 92134 32048 92218
rect 31728 91898 31770 92134
rect 32006 91898 32048 92134
rect 31728 91876 32048 91898
rect 62448 92454 62768 92476
rect 62448 92218 62490 92454
rect 62726 92218 62768 92454
rect 62448 92134 62768 92218
rect 62448 91898 62490 92134
rect 62726 91898 62768 92134
rect 62448 91876 62768 91898
rect 93168 92454 93488 92476
rect 93168 92218 93210 92454
rect 93446 92218 93488 92454
rect 93168 92134 93488 92218
rect 93168 91898 93210 92134
rect 93446 91898 93488 92134
rect 93168 91876 93488 91898
rect 123888 92454 124208 92476
rect 123888 92218 123930 92454
rect 124166 92218 124208 92454
rect 123888 92134 124208 92218
rect 123888 91898 123930 92134
rect 124166 91898 124208 92134
rect 123888 91876 124208 91898
rect 154608 92454 154928 92476
rect 154608 92218 154650 92454
rect 154886 92218 154928 92454
rect 154608 92134 154928 92218
rect 154608 91898 154650 92134
rect 154886 91898 154928 92134
rect 154608 91876 154928 91898
rect 185328 92454 185648 92476
rect 185328 92218 185370 92454
rect 185606 92218 185648 92454
rect 185328 92134 185648 92218
rect 185328 91898 185370 92134
rect 185606 91898 185648 92134
rect 185328 91876 185648 91898
rect 216048 92454 216368 92476
rect 216048 92218 216090 92454
rect 216326 92218 216368 92454
rect 216048 92134 216368 92218
rect 216048 91898 216090 92134
rect 216326 91898 216368 92134
rect 216048 91876 216368 91898
rect 246768 92454 247088 92476
rect 246768 92218 246810 92454
rect 247046 92218 247088 92454
rect 246768 92134 247088 92218
rect 246768 91898 246810 92134
rect 247046 91898 247088 92134
rect 246768 91876 247088 91898
rect 270804 92454 271404 127898
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1286 19404 19898
rect 18804 -1522 18986 -1286
rect 19222 -1522 19404 -1286
rect 18804 -1606 19404 -1522
rect 18804 -1842 18986 -1606
rect 19222 -1842 19404 -1606
rect 18804 -1864 19404 -1842
rect 36804 38454 37404 72600
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1864 37404 -902
rect 54804 56454 55404 72600
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1286 55404 19898
rect 54804 -1522 54986 -1286
rect 55222 -1522 55404 -1286
rect 54804 -1606 55404 -1522
rect 54804 -1842 54986 -1606
rect 55222 -1842 55404 -1606
rect 54804 -1864 55404 -1842
rect 72804 38454 73404 72600
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1864 73404 -902
rect 90804 56454 91404 72600
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1286 91404 19898
rect 90804 -1522 90986 -1286
rect 91222 -1522 91404 -1286
rect 90804 -1606 91404 -1522
rect 90804 -1842 90986 -1606
rect 91222 -1842 91404 -1606
rect 90804 -1864 91404 -1842
rect 108804 38454 109404 72600
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1864 109404 -902
rect 126804 56454 127404 72600
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1286 127404 19898
rect 126804 -1522 126986 -1286
rect 127222 -1522 127404 -1286
rect 126804 -1606 127404 -1522
rect 126804 -1842 126986 -1606
rect 127222 -1842 127404 -1606
rect 126804 -1864 127404 -1842
rect 144804 38454 145404 72600
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1864 145404 -902
rect 162804 56454 163404 72600
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1286 163404 19898
rect 162804 -1522 162986 -1286
rect 163222 -1522 163404 -1286
rect 162804 -1606 163404 -1522
rect 162804 -1842 162986 -1606
rect 163222 -1842 163404 -1606
rect 162804 -1864 163404 -1842
rect 180804 38454 181404 72600
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1864 181404 -902
rect 198804 56454 199404 72600
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1286 199404 19898
rect 198804 -1522 198986 -1286
rect 199222 -1522 199404 -1286
rect 198804 -1606 199404 -1522
rect 198804 -1842 198986 -1606
rect 199222 -1842 199404 -1606
rect 198804 -1864 199404 -1842
rect 216804 38454 217404 72600
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1864 217404 -902
rect 234804 56454 235404 72600
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 234804 20454 235404 55898
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1286 235404 19898
rect 234804 -1522 234986 -1286
rect 235222 -1522 235404 -1286
rect 234804 -1606 235404 -1522
rect 234804 -1842 234986 -1606
rect 235222 -1842 235404 -1606
rect 234804 -1864 235404 -1842
rect 252804 38454 253404 72600
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1864 253404 -902
rect 270804 56454 271404 91898
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1286 271404 19898
rect 270804 -1522 270986 -1286
rect 271222 -1522 271404 -1286
rect 270804 -1606 271404 -1522
rect 270804 -1842 270986 -1606
rect 271222 -1842 271404 -1606
rect 270804 -1864 271404 -1842
rect 288804 290454 289404 314560
rect 288804 290218 288986 290454
rect 289222 290218 289404 290454
rect 288804 290134 289404 290218
rect 288804 289898 288986 290134
rect 289222 289898 289404 290134
rect 288804 254454 289404 289898
rect 288804 254218 288986 254454
rect 289222 254218 289404 254454
rect 288804 254134 289404 254218
rect 288804 253898 288986 254134
rect 289222 253898 289404 254134
rect 288804 218454 289404 253898
rect 288804 218218 288986 218454
rect 289222 218218 289404 218454
rect 288804 218134 289404 218218
rect 288804 217898 288986 218134
rect 289222 217898 289404 218134
rect 288804 182454 289404 217898
rect 288804 182218 288986 182454
rect 289222 182218 289404 182454
rect 288804 182134 289404 182218
rect 288804 181898 288986 182134
rect 289222 181898 289404 182134
rect 288804 146454 289404 181898
rect 288804 146218 288986 146454
rect 289222 146218 289404 146454
rect 288804 146134 289404 146218
rect 288804 145898 288986 146134
rect 289222 145898 289404 146134
rect 288804 110454 289404 145898
rect 288804 110218 288986 110454
rect 289222 110218 289404 110454
rect 288804 110134 289404 110218
rect 288804 109898 288986 110134
rect 289222 109898 289404 110134
rect 288804 74454 289404 109898
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 288804 38454 289404 73898
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1864 289404 -902
rect 306804 308454 307404 314560
rect 306804 308218 306986 308454
rect 307222 308218 307404 308454
rect 306804 308134 307404 308218
rect 306804 307898 306986 308134
rect 307222 307898 307404 308134
rect 306804 272454 307404 307898
rect 324804 290454 325404 325898
rect 324804 290218 324986 290454
rect 325222 290218 325404 290454
rect 324804 290134 325404 290218
rect 324804 289898 324986 290134
rect 325222 289898 325404 290134
rect 324804 274600 325404 289898
rect 342804 380454 343404 382916
rect 342804 380218 342986 380454
rect 343222 380218 343404 380454
rect 342804 380134 343404 380218
rect 342804 379898 342986 380134
rect 343222 379898 343404 380134
rect 342804 344454 343404 379898
rect 342804 344218 342986 344454
rect 343222 344218 343404 344454
rect 342804 344134 343404 344218
rect 342804 343898 342986 344134
rect 343222 343898 343404 344134
rect 342804 308454 343404 343898
rect 342804 308218 342986 308454
rect 343222 308218 343404 308454
rect 342804 308134 343404 308218
rect 342804 307898 342986 308134
rect 343222 307898 343404 308134
rect 342804 274600 343404 307898
rect 360804 362454 361404 382916
rect 360804 362218 360986 362454
rect 361222 362218 361404 362454
rect 360804 362134 361404 362218
rect 360804 361898 360986 362134
rect 361222 361898 361404 362134
rect 360804 326454 361404 361898
rect 360804 326218 360986 326454
rect 361222 326218 361404 326454
rect 360804 326134 361404 326218
rect 360804 325898 360986 326134
rect 361222 325898 361404 326134
rect 360804 290454 361404 325898
rect 360804 290218 360986 290454
rect 361222 290218 361404 290454
rect 360804 290134 361404 290218
rect 360804 289898 360986 290134
rect 361222 289898 361404 290134
rect 360804 274600 361404 289898
rect 378804 380454 379404 382916
rect 378804 380218 378986 380454
rect 379222 380218 379404 380454
rect 378804 380134 379404 380218
rect 378804 379898 378986 380134
rect 379222 379898 379404 380134
rect 378804 344454 379404 379898
rect 378804 344218 378986 344454
rect 379222 344218 379404 344454
rect 378804 344134 379404 344218
rect 378804 343898 378986 344134
rect 379222 343898 379404 344134
rect 378804 308454 379404 343898
rect 378804 308218 378986 308454
rect 379222 308218 379404 308454
rect 378804 308134 379404 308218
rect 378804 307898 378986 308134
rect 379222 307898 379404 308134
rect 378804 274600 379404 307898
rect 396804 362454 397404 382916
rect 396804 362218 396986 362454
rect 397222 362218 397404 362454
rect 396804 362134 397404 362218
rect 396804 361898 396986 362134
rect 397222 361898 397404 362134
rect 396804 326454 397404 361898
rect 396804 326218 396986 326454
rect 397222 326218 397404 326454
rect 396804 326134 397404 326218
rect 396804 325898 396986 326134
rect 397222 325898 397404 326134
rect 396804 290454 397404 325898
rect 396804 290218 396986 290454
rect 397222 290218 397404 290454
rect 396804 290134 397404 290218
rect 396804 289898 396986 290134
rect 397222 289898 397404 290134
rect 396804 274600 397404 289898
rect 414804 380454 415404 382916
rect 414804 380218 414986 380454
rect 415222 380218 415404 380454
rect 414804 380134 415404 380218
rect 414804 379898 414986 380134
rect 415222 379898 415404 380134
rect 414804 344454 415404 379898
rect 414804 344218 414986 344454
rect 415222 344218 415404 344454
rect 414804 344134 415404 344218
rect 414804 343898 414986 344134
rect 415222 343898 415404 344134
rect 414804 308454 415404 343898
rect 414804 308218 414986 308454
rect 415222 308218 415404 308454
rect 414804 308134 415404 308218
rect 414804 307898 414986 308134
rect 415222 307898 415404 308134
rect 414804 274600 415404 307898
rect 432804 362454 433404 382916
rect 432804 362218 432986 362454
rect 433222 362218 433404 362454
rect 432804 362134 433404 362218
rect 432804 361898 432986 362134
rect 433222 361898 433404 362134
rect 432804 326454 433404 361898
rect 432804 326218 432986 326454
rect 433222 326218 433404 326454
rect 432804 326134 433404 326218
rect 432804 325898 432986 326134
rect 433222 325898 433404 326134
rect 432804 290454 433404 325898
rect 432804 290218 432986 290454
rect 433222 290218 433404 290454
rect 432804 290134 433404 290218
rect 432804 289898 432986 290134
rect 433222 289898 433404 290134
rect 432804 274600 433404 289898
rect 450804 380454 451404 382916
rect 450804 380218 450986 380454
rect 451222 380218 451404 380454
rect 450804 380134 451404 380218
rect 450804 379898 450986 380134
rect 451222 379898 451404 380134
rect 450804 344454 451404 379898
rect 450804 344218 450986 344454
rect 451222 344218 451404 344454
rect 450804 344134 451404 344218
rect 450804 343898 450986 344134
rect 451222 343898 451404 344134
rect 450804 308454 451404 343898
rect 450804 308218 450986 308454
rect 451222 308218 451404 308454
rect 450804 308134 451404 308218
rect 450804 307898 450986 308134
rect 451222 307898 451404 308134
rect 450804 274600 451404 307898
rect 468804 362454 469404 382916
rect 468804 362218 468986 362454
rect 469222 362218 469404 362454
rect 468804 362134 469404 362218
rect 468804 361898 468986 362134
rect 469222 361898 469404 362134
rect 468804 326454 469404 361898
rect 468804 326218 468986 326454
rect 469222 326218 469404 326454
rect 468804 326134 469404 326218
rect 468804 325898 468986 326134
rect 469222 325898 469404 326134
rect 468804 290454 469404 325898
rect 468804 290218 468986 290454
rect 469222 290218 469404 290454
rect 468804 290134 469404 290218
rect 468804 289898 468986 290134
rect 469222 289898 469404 290134
rect 468804 274600 469404 289898
rect 486804 380454 487404 382916
rect 486804 380218 486986 380454
rect 487222 380218 487404 380454
rect 486804 380134 487404 380218
rect 486804 379898 486986 380134
rect 487222 379898 487404 380134
rect 486804 344454 487404 379898
rect 486804 344218 486986 344454
rect 487222 344218 487404 344454
rect 486804 344134 487404 344218
rect 486804 343898 486986 344134
rect 487222 343898 487404 344134
rect 486804 308454 487404 343898
rect 486804 308218 486986 308454
rect 487222 308218 487404 308454
rect 486804 308134 487404 308218
rect 486804 307898 486986 308134
rect 487222 307898 487404 308134
rect 486804 274600 487404 307898
rect 504804 362454 505404 382916
rect 504804 362218 504986 362454
rect 505222 362218 505404 362454
rect 504804 362134 505404 362218
rect 504804 361898 504986 362134
rect 505222 361898 505404 362134
rect 504804 326454 505404 361898
rect 504804 326218 504986 326454
rect 505222 326218 505404 326454
rect 504804 326134 505404 326218
rect 504804 325898 504986 326134
rect 505222 325898 505404 326134
rect 504804 290454 505404 325898
rect 504804 290218 504986 290454
rect 505222 290218 505404 290454
rect 504804 290134 505404 290218
rect 504804 289898 504986 290134
rect 505222 289898 505404 290134
rect 504804 274600 505404 289898
rect 522804 380454 523404 382916
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 274600 523404 307898
rect 540804 362454 541404 382916
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 274600 541404 289898
rect 558804 380454 559404 382916
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 274600 559404 307898
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 306804 272218 306986 272454
rect 307222 272218 307404 272454
rect 306804 272134 307404 272218
rect 306804 271898 306986 272134
rect 307222 271898 307404 272134
rect 306804 236454 307404 271898
rect 339216 254454 339536 254476
rect 339216 254218 339258 254454
rect 339494 254218 339536 254454
rect 339216 254134 339536 254218
rect 339216 253898 339258 254134
rect 339494 253898 339536 254134
rect 339216 253876 339536 253898
rect 369936 254454 370256 254476
rect 369936 254218 369978 254454
rect 370214 254218 370256 254454
rect 369936 254134 370256 254218
rect 369936 253898 369978 254134
rect 370214 253898 370256 254134
rect 369936 253876 370256 253898
rect 400656 254454 400976 254476
rect 400656 254218 400698 254454
rect 400934 254218 400976 254454
rect 400656 254134 400976 254218
rect 400656 253898 400698 254134
rect 400934 253898 400976 254134
rect 400656 253876 400976 253898
rect 431376 254454 431696 254476
rect 431376 254218 431418 254454
rect 431654 254218 431696 254454
rect 431376 254134 431696 254218
rect 431376 253898 431418 254134
rect 431654 253898 431696 254134
rect 431376 253876 431696 253898
rect 462096 254454 462416 254476
rect 462096 254218 462138 254454
rect 462374 254218 462416 254454
rect 462096 254134 462416 254218
rect 462096 253898 462138 254134
rect 462374 253898 462416 254134
rect 462096 253876 462416 253898
rect 492816 254454 493136 254476
rect 492816 254218 492858 254454
rect 493094 254218 493136 254454
rect 492816 254134 493136 254218
rect 492816 253898 492858 254134
rect 493094 253898 493136 254134
rect 492816 253876 493136 253898
rect 523536 254454 523856 254476
rect 523536 254218 523578 254454
rect 523814 254218 523856 254454
rect 523536 254134 523856 254218
rect 523536 253898 523578 254134
rect 523814 253898 523856 254134
rect 523536 253876 523856 253898
rect 554256 254454 554576 254476
rect 554256 254218 554298 254454
rect 554534 254218 554576 254454
rect 554256 254134 554576 254218
rect 554256 253898 554298 254134
rect 554534 253898 554576 254134
rect 554256 253876 554576 253898
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 306804 236218 306986 236454
rect 307222 236218 307404 236454
rect 306804 236134 307404 236218
rect 306804 235898 306986 236134
rect 307222 235898 307404 236134
rect 306804 200454 307404 235898
rect 323856 236454 324176 236476
rect 323856 236218 323898 236454
rect 324134 236218 324176 236454
rect 323856 236134 324176 236218
rect 323856 235898 323898 236134
rect 324134 235898 324176 236134
rect 323856 235876 324176 235898
rect 354576 236454 354896 236476
rect 354576 236218 354618 236454
rect 354854 236218 354896 236454
rect 354576 236134 354896 236218
rect 354576 235898 354618 236134
rect 354854 235898 354896 236134
rect 354576 235876 354896 235898
rect 385296 236454 385616 236476
rect 385296 236218 385338 236454
rect 385574 236218 385616 236454
rect 385296 236134 385616 236218
rect 385296 235898 385338 236134
rect 385574 235898 385616 236134
rect 385296 235876 385616 235898
rect 416016 236454 416336 236476
rect 416016 236218 416058 236454
rect 416294 236218 416336 236454
rect 416016 236134 416336 236218
rect 416016 235898 416058 236134
rect 416294 235898 416336 236134
rect 416016 235876 416336 235898
rect 446736 236454 447056 236476
rect 446736 236218 446778 236454
rect 447014 236218 447056 236454
rect 446736 236134 447056 236218
rect 446736 235898 446778 236134
rect 447014 235898 447056 236134
rect 446736 235876 447056 235898
rect 477456 236454 477776 236476
rect 477456 236218 477498 236454
rect 477734 236218 477776 236454
rect 477456 236134 477776 236218
rect 477456 235898 477498 236134
rect 477734 235898 477776 236134
rect 477456 235876 477776 235898
rect 508176 236454 508496 236476
rect 508176 236218 508218 236454
rect 508454 236218 508496 236454
rect 508176 236134 508496 236218
rect 508176 235898 508218 236134
rect 508454 235898 508496 236134
rect 508176 235876 508496 235898
rect 538896 236454 539216 236476
rect 538896 236218 538938 236454
rect 539174 236218 539216 236454
rect 538896 236134 539216 236218
rect 538896 235898 538938 236134
rect 539174 235898 539216 236134
rect 538896 235876 539216 235898
rect 339216 218454 339536 218476
rect 339216 218218 339258 218454
rect 339494 218218 339536 218454
rect 339216 218134 339536 218218
rect 339216 217898 339258 218134
rect 339494 217898 339536 218134
rect 339216 217876 339536 217898
rect 369936 218454 370256 218476
rect 369936 218218 369978 218454
rect 370214 218218 370256 218454
rect 369936 218134 370256 218218
rect 369936 217898 369978 218134
rect 370214 217898 370256 218134
rect 369936 217876 370256 217898
rect 400656 218454 400976 218476
rect 400656 218218 400698 218454
rect 400934 218218 400976 218454
rect 400656 218134 400976 218218
rect 400656 217898 400698 218134
rect 400934 217898 400976 218134
rect 400656 217876 400976 217898
rect 431376 218454 431696 218476
rect 431376 218218 431418 218454
rect 431654 218218 431696 218454
rect 431376 218134 431696 218218
rect 431376 217898 431418 218134
rect 431654 217898 431696 218134
rect 431376 217876 431696 217898
rect 462096 218454 462416 218476
rect 462096 218218 462138 218454
rect 462374 218218 462416 218454
rect 462096 218134 462416 218218
rect 462096 217898 462138 218134
rect 462374 217898 462416 218134
rect 462096 217876 462416 217898
rect 492816 218454 493136 218476
rect 492816 218218 492858 218454
rect 493094 218218 493136 218454
rect 492816 218134 493136 218218
rect 492816 217898 492858 218134
rect 493094 217898 493136 218134
rect 492816 217876 493136 217898
rect 523536 218454 523856 218476
rect 523536 218218 523578 218454
rect 523814 218218 523856 218454
rect 523536 218134 523856 218218
rect 523536 217898 523578 218134
rect 523814 217898 523856 218134
rect 523536 217876 523856 217898
rect 554256 218454 554576 218476
rect 554256 218218 554298 218454
rect 554534 218218 554576 218454
rect 554256 218134 554576 218218
rect 554256 217898 554298 218134
rect 554534 217898 554576 218134
rect 554256 217876 554576 217898
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 306804 200218 306986 200454
rect 307222 200218 307404 200454
rect 306804 200134 307404 200218
rect 306804 199898 306986 200134
rect 307222 199898 307404 200134
rect 306804 164454 307404 199898
rect 323856 200454 324176 200476
rect 323856 200218 323898 200454
rect 324134 200218 324176 200454
rect 323856 200134 324176 200218
rect 323856 199898 323898 200134
rect 324134 199898 324176 200134
rect 323856 199876 324176 199898
rect 354576 200454 354896 200476
rect 354576 200218 354618 200454
rect 354854 200218 354896 200454
rect 354576 200134 354896 200218
rect 354576 199898 354618 200134
rect 354854 199898 354896 200134
rect 354576 199876 354896 199898
rect 385296 200454 385616 200476
rect 385296 200218 385338 200454
rect 385574 200218 385616 200454
rect 385296 200134 385616 200218
rect 385296 199898 385338 200134
rect 385574 199898 385616 200134
rect 385296 199876 385616 199898
rect 416016 200454 416336 200476
rect 416016 200218 416058 200454
rect 416294 200218 416336 200454
rect 416016 200134 416336 200218
rect 416016 199898 416058 200134
rect 416294 199898 416336 200134
rect 416016 199876 416336 199898
rect 446736 200454 447056 200476
rect 446736 200218 446778 200454
rect 447014 200218 447056 200454
rect 446736 200134 447056 200218
rect 446736 199898 446778 200134
rect 447014 199898 447056 200134
rect 446736 199876 447056 199898
rect 477456 200454 477776 200476
rect 477456 200218 477498 200454
rect 477734 200218 477776 200454
rect 477456 200134 477776 200218
rect 477456 199898 477498 200134
rect 477734 199898 477776 200134
rect 477456 199876 477776 199898
rect 508176 200454 508496 200476
rect 508176 200218 508218 200454
rect 508454 200218 508496 200454
rect 508176 200134 508496 200218
rect 508176 199898 508218 200134
rect 508454 199898 508496 200134
rect 508176 199876 508496 199898
rect 538896 200454 539216 200476
rect 538896 200218 538938 200454
rect 539174 200218 539216 200454
rect 538896 200134 539216 200218
rect 538896 199898 538938 200134
rect 539174 199898 539216 200134
rect 538896 199876 539216 199898
rect 339216 182454 339536 182476
rect 339216 182218 339258 182454
rect 339494 182218 339536 182454
rect 339216 182134 339536 182218
rect 339216 181898 339258 182134
rect 339494 181898 339536 182134
rect 339216 181876 339536 181898
rect 369936 182454 370256 182476
rect 369936 182218 369978 182454
rect 370214 182218 370256 182454
rect 369936 182134 370256 182218
rect 369936 181898 369978 182134
rect 370214 181898 370256 182134
rect 369936 181876 370256 181898
rect 400656 182454 400976 182476
rect 400656 182218 400698 182454
rect 400934 182218 400976 182454
rect 400656 182134 400976 182218
rect 400656 181898 400698 182134
rect 400934 181898 400976 182134
rect 400656 181876 400976 181898
rect 431376 182454 431696 182476
rect 431376 182218 431418 182454
rect 431654 182218 431696 182454
rect 431376 182134 431696 182218
rect 431376 181898 431418 182134
rect 431654 181898 431696 182134
rect 431376 181876 431696 181898
rect 462096 182454 462416 182476
rect 462096 182218 462138 182454
rect 462374 182218 462416 182454
rect 462096 182134 462416 182218
rect 462096 181898 462138 182134
rect 462374 181898 462416 182134
rect 462096 181876 462416 181898
rect 492816 182454 493136 182476
rect 492816 182218 492858 182454
rect 493094 182218 493136 182454
rect 492816 182134 493136 182218
rect 492816 181898 492858 182134
rect 493094 181898 493136 182134
rect 492816 181876 493136 181898
rect 523536 182454 523856 182476
rect 523536 182218 523578 182454
rect 523814 182218 523856 182454
rect 523536 182134 523856 182218
rect 523536 181898 523578 182134
rect 523814 181898 523856 182134
rect 523536 181876 523856 181898
rect 554256 182454 554576 182476
rect 554256 182218 554298 182454
rect 554534 182218 554576 182454
rect 554256 182134 554576 182218
rect 554256 181898 554298 182134
rect 554534 181898 554576 182134
rect 554256 181876 554576 181898
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 306804 164218 306986 164454
rect 307222 164218 307404 164454
rect 306804 164134 307404 164218
rect 306804 163898 306986 164134
rect 307222 163898 307404 164134
rect 306804 128454 307404 163898
rect 323856 164454 324176 164476
rect 323856 164218 323898 164454
rect 324134 164218 324176 164454
rect 323856 164134 324176 164218
rect 323856 163898 323898 164134
rect 324134 163898 324176 164134
rect 323856 163876 324176 163898
rect 354576 164454 354896 164476
rect 354576 164218 354618 164454
rect 354854 164218 354896 164454
rect 354576 164134 354896 164218
rect 354576 163898 354618 164134
rect 354854 163898 354896 164134
rect 354576 163876 354896 163898
rect 385296 164454 385616 164476
rect 385296 164218 385338 164454
rect 385574 164218 385616 164454
rect 385296 164134 385616 164218
rect 385296 163898 385338 164134
rect 385574 163898 385616 164134
rect 385296 163876 385616 163898
rect 416016 164454 416336 164476
rect 416016 164218 416058 164454
rect 416294 164218 416336 164454
rect 416016 164134 416336 164218
rect 416016 163898 416058 164134
rect 416294 163898 416336 164134
rect 416016 163876 416336 163898
rect 446736 164454 447056 164476
rect 446736 164218 446778 164454
rect 447014 164218 447056 164454
rect 446736 164134 447056 164218
rect 446736 163898 446778 164134
rect 447014 163898 447056 164134
rect 446736 163876 447056 163898
rect 477456 164454 477776 164476
rect 477456 164218 477498 164454
rect 477734 164218 477776 164454
rect 477456 164134 477776 164218
rect 477456 163898 477498 164134
rect 477734 163898 477776 164134
rect 477456 163876 477776 163898
rect 508176 164454 508496 164476
rect 508176 164218 508218 164454
rect 508454 164218 508496 164454
rect 508176 164134 508496 164218
rect 508176 163898 508218 164134
rect 508454 163898 508496 164134
rect 508176 163876 508496 163898
rect 538896 164454 539216 164476
rect 538896 164218 538938 164454
rect 539174 164218 539216 164454
rect 538896 164134 539216 164218
rect 538896 163898 538938 164134
rect 539174 163898 539216 164134
rect 538896 163876 539216 163898
rect 339216 146454 339536 146476
rect 339216 146218 339258 146454
rect 339494 146218 339536 146454
rect 339216 146134 339536 146218
rect 339216 145898 339258 146134
rect 339494 145898 339536 146134
rect 339216 145876 339536 145898
rect 369936 146454 370256 146476
rect 369936 146218 369978 146454
rect 370214 146218 370256 146454
rect 369936 146134 370256 146218
rect 369936 145898 369978 146134
rect 370214 145898 370256 146134
rect 369936 145876 370256 145898
rect 400656 146454 400976 146476
rect 400656 146218 400698 146454
rect 400934 146218 400976 146454
rect 400656 146134 400976 146218
rect 400656 145898 400698 146134
rect 400934 145898 400976 146134
rect 400656 145876 400976 145898
rect 431376 146454 431696 146476
rect 431376 146218 431418 146454
rect 431654 146218 431696 146454
rect 431376 146134 431696 146218
rect 431376 145898 431418 146134
rect 431654 145898 431696 146134
rect 431376 145876 431696 145898
rect 462096 146454 462416 146476
rect 462096 146218 462138 146454
rect 462374 146218 462416 146454
rect 462096 146134 462416 146218
rect 462096 145898 462138 146134
rect 462374 145898 462416 146134
rect 462096 145876 462416 145898
rect 492816 146454 493136 146476
rect 492816 146218 492858 146454
rect 493094 146218 493136 146454
rect 492816 146134 493136 146218
rect 492816 145898 492858 146134
rect 493094 145898 493136 146134
rect 492816 145876 493136 145898
rect 523536 146454 523856 146476
rect 523536 146218 523578 146454
rect 523814 146218 523856 146454
rect 523536 146134 523856 146218
rect 523536 145898 523578 146134
rect 523814 145898 523856 146134
rect 523536 145876 523856 145898
rect 554256 146454 554576 146476
rect 554256 146218 554298 146454
rect 554534 146218 554576 146454
rect 554256 146134 554576 146218
rect 554256 145898 554298 146134
rect 554534 145898 554576 146134
rect 554256 145876 554576 145898
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 306804 128218 306986 128454
rect 307222 128218 307404 128454
rect 306804 128134 307404 128218
rect 306804 127898 306986 128134
rect 307222 127898 307404 128134
rect 306804 92454 307404 127898
rect 323856 128454 324176 128476
rect 323856 128218 323898 128454
rect 324134 128218 324176 128454
rect 323856 128134 324176 128218
rect 323856 127898 323898 128134
rect 324134 127898 324176 128134
rect 323856 127876 324176 127898
rect 354576 128454 354896 128476
rect 354576 128218 354618 128454
rect 354854 128218 354896 128454
rect 354576 128134 354896 128218
rect 354576 127898 354618 128134
rect 354854 127898 354896 128134
rect 354576 127876 354896 127898
rect 385296 128454 385616 128476
rect 385296 128218 385338 128454
rect 385574 128218 385616 128454
rect 385296 128134 385616 128218
rect 385296 127898 385338 128134
rect 385574 127898 385616 128134
rect 385296 127876 385616 127898
rect 416016 128454 416336 128476
rect 416016 128218 416058 128454
rect 416294 128218 416336 128454
rect 416016 128134 416336 128218
rect 416016 127898 416058 128134
rect 416294 127898 416336 128134
rect 416016 127876 416336 127898
rect 446736 128454 447056 128476
rect 446736 128218 446778 128454
rect 447014 128218 447056 128454
rect 446736 128134 447056 128218
rect 446736 127898 446778 128134
rect 447014 127898 447056 128134
rect 446736 127876 447056 127898
rect 477456 128454 477776 128476
rect 477456 128218 477498 128454
rect 477734 128218 477776 128454
rect 477456 128134 477776 128218
rect 477456 127898 477498 128134
rect 477734 127898 477776 128134
rect 477456 127876 477776 127898
rect 508176 128454 508496 128476
rect 508176 128218 508218 128454
rect 508454 128218 508496 128454
rect 508176 128134 508496 128218
rect 508176 127898 508218 128134
rect 508454 127898 508496 128134
rect 508176 127876 508496 127898
rect 538896 128454 539216 128476
rect 538896 128218 538938 128454
rect 539174 128218 539216 128454
rect 538896 128134 539216 128218
rect 538896 127898 538938 128134
rect 539174 127898 539216 128134
rect 538896 127876 539216 127898
rect 339216 110454 339536 110476
rect 339216 110218 339258 110454
rect 339494 110218 339536 110454
rect 339216 110134 339536 110218
rect 339216 109898 339258 110134
rect 339494 109898 339536 110134
rect 339216 109876 339536 109898
rect 369936 110454 370256 110476
rect 369936 110218 369978 110454
rect 370214 110218 370256 110454
rect 369936 110134 370256 110218
rect 369936 109898 369978 110134
rect 370214 109898 370256 110134
rect 369936 109876 370256 109898
rect 400656 110454 400976 110476
rect 400656 110218 400698 110454
rect 400934 110218 400976 110454
rect 400656 110134 400976 110218
rect 400656 109898 400698 110134
rect 400934 109898 400976 110134
rect 400656 109876 400976 109898
rect 431376 110454 431696 110476
rect 431376 110218 431418 110454
rect 431654 110218 431696 110454
rect 431376 110134 431696 110218
rect 431376 109898 431418 110134
rect 431654 109898 431696 110134
rect 431376 109876 431696 109898
rect 462096 110454 462416 110476
rect 462096 110218 462138 110454
rect 462374 110218 462416 110454
rect 462096 110134 462416 110218
rect 462096 109898 462138 110134
rect 462374 109898 462416 110134
rect 462096 109876 462416 109898
rect 492816 110454 493136 110476
rect 492816 110218 492858 110454
rect 493094 110218 493136 110454
rect 492816 110134 493136 110218
rect 492816 109898 492858 110134
rect 493094 109898 493136 110134
rect 492816 109876 493136 109898
rect 523536 110454 523856 110476
rect 523536 110218 523578 110454
rect 523814 110218 523856 110454
rect 523536 110134 523856 110218
rect 523536 109898 523578 110134
rect 523814 109898 523856 110134
rect 523536 109876 523856 109898
rect 554256 110454 554576 110476
rect 554256 110218 554298 110454
rect 554534 110218 554576 110454
rect 554256 110134 554576 110218
rect 554256 109898 554298 110134
rect 554534 109898 554576 110134
rect 554256 109876 554576 109898
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 306804 56454 307404 91898
rect 323856 92454 324176 92476
rect 323856 92218 323898 92454
rect 324134 92218 324176 92454
rect 323856 92134 324176 92218
rect 323856 91898 323898 92134
rect 324134 91898 324176 92134
rect 323856 91876 324176 91898
rect 354576 92454 354896 92476
rect 354576 92218 354618 92454
rect 354854 92218 354896 92454
rect 354576 92134 354896 92218
rect 354576 91898 354618 92134
rect 354854 91898 354896 92134
rect 354576 91876 354896 91898
rect 385296 92454 385616 92476
rect 385296 92218 385338 92454
rect 385574 92218 385616 92454
rect 385296 92134 385616 92218
rect 385296 91898 385338 92134
rect 385574 91898 385616 92134
rect 385296 91876 385616 91898
rect 416016 92454 416336 92476
rect 416016 92218 416058 92454
rect 416294 92218 416336 92454
rect 416016 92134 416336 92218
rect 416016 91898 416058 92134
rect 416294 91898 416336 92134
rect 416016 91876 416336 91898
rect 446736 92454 447056 92476
rect 446736 92218 446778 92454
rect 447014 92218 447056 92454
rect 446736 92134 447056 92218
rect 446736 91898 446778 92134
rect 447014 91898 447056 92134
rect 446736 91876 447056 91898
rect 477456 92454 477776 92476
rect 477456 92218 477498 92454
rect 477734 92218 477776 92454
rect 477456 92134 477776 92218
rect 477456 91898 477498 92134
rect 477734 91898 477776 92134
rect 477456 91876 477776 91898
rect 508176 92454 508496 92476
rect 508176 92218 508218 92454
rect 508454 92218 508496 92454
rect 508176 92134 508496 92218
rect 508176 91898 508218 92134
rect 508454 91898 508496 92134
rect 508176 91876 508496 91898
rect 538896 92454 539216 92476
rect 538896 92218 538938 92454
rect 539174 92218 539216 92454
rect 538896 92134 539216 92218
rect 538896 91898 538938 92134
rect 539174 91898 539216 92134
rect 538896 91876 539216 91898
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1286 307404 19898
rect 306804 -1522 306986 -1286
rect 307222 -1522 307404 -1286
rect 306804 -1606 307404 -1522
rect 306804 -1842 306986 -1606
rect 307222 -1842 307404 -1606
rect 306804 -1864 307404 -1842
rect 324804 38454 325404 72600
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1864 325404 -902
rect 342804 56454 343404 72600
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1286 343404 19898
rect 342804 -1522 342986 -1286
rect 343222 -1522 343404 -1286
rect 342804 -1606 343404 -1522
rect 342804 -1842 342986 -1606
rect 343222 -1842 343404 -1606
rect 342804 -1864 343404 -1842
rect 360804 38454 361404 72600
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1864 361404 -902
rect 378804 56454 379404 72600
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1286 379404 19898
rect 378804 -1522 378986 -1286
rect 379222 -1522 379404 -1286
rect 378804 -1606 379404 -1522
rect 378804 -1842 378986 -1606
rect 379222 -1842 379404 -1606
rect 378804 -1864 379404 -1842
rect 396804 38454 397404 72600
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1864 397404 -902
rect 414804 56454 415404 72600
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1286 415404 19898
rect 414804 -1522 414986 -1286
rect 415222 -1522 415404 -1286
rect 414804 -1606 415404 -1522
rect 414804 -1842 414986 -1606
rect 415222 -1842 415404 -1606
rect 414804 -1864 415404 -1842
rect 432804 38454 433404 72600
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1864 433404 -902
rect 450804 56454 451404 72600
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1286 451404 19898
rect 450804 -1522 450986 -1286
rect 451222 -1522 451404 -1286
rect 450804 -1606 451404 -1522
rect 450804 -1842 450986 -1606
rect 451222 -1842 451404 -1606
rect 450804 -1864 451404 -1842
rect 468804 38454 469404 72600
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1864 469404 -902
rect 486804 56454 487404 72600
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1286 487404 19898
rect 486804 -1522 486986 -1286
rect 487222 -1522 487404 -1286
rect 486804 -1606 487404 -1522
rect 486804 -1842 486986 -1606
rect 487222 -1842 487404 -1606
rect 486804 -1864 487404 -1842
rect 504804 38454 505404 72600
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1864 505404 -902
rect 522804 56454 523404 72600
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1286 523404 19898
rect 522804 -1522 522986 -1286
rect 523222 -1522 523404 -1286
rect 522804 -1606 523404 -1522
rect 522804 -1842 522986 -1606
rect 523222 -1842 523404 -1606
rect 522804 -1864 523404 -1842
rect 540804 38454 541404 72600
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1864 541404 -902
rect 558804 56454 559404 72600
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1286 559404 19898
rect 558804 -1522 558986 -1286
rect 559222 -1522 559404 -1286
rect 558804 -1606 559404 -1522
rect 558804 -1842 558986 -1606
rect 559222 -1842 559404 -1606
rect 558804 -1864 559404 -1842
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1864 577404 -902
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586260 668454 586860 705222
rect 586260 668218 586442 668454
rect 586678 668218 586860 668454
rect 586260 668134 586860 668218
rect 586260 667898 586442 668134
rect 586678 667898 586860 668134
rect 586260 632454 586860 667898
rect 586260 632218 586442 632454
rect 586678 632218 586860 632454
rect 586260 632134 586860 632218
rect 586260 631898 586442 632134
rect 586678 631898 586860 632134
rect 586260 596454 586860 631898
rect 586260 596218 586442 596454
rect 586678 596218 586860 596454
rect 586260 596134 586860 596218
rect 586260 595898 586442 596134
rect 586678 595898 586860 596134
rect 586260 560454 586860 595898
rect 586260 560218 586442 560454
rect 586678 560218 586860 560454
rect 586260 560134 586860 560218
rect 586260 559898 586442 560134
rect 586678 559898 586860 560134
rect 586260 524454 586860 559898
rect 586260 524218 586442 524454
rect 586678 524218 586860 524454
rect 586260 524134 586860 524218
rect 586260 523898 586442 524134
rect 586678 523898 586860 524134
rect 586260 488454 586860 523898
rect 586260 488218 586442 488454
rect 586678 488218 586860 488454
rect 586260 488134 586860 488218
rect 586260 487898 586442 488134
rect 586678 487898 586860 488134
rect 586260 452454 586860 487898
rect 586260 452218 586442 452454
rect 586678 452218 586860 452454
rect 586260 452134 586860 452218
rect 586260 451898 586442 452134
rect 586678 451898 586860 452134
rect 586260 416454 586860 451898
rect 586260 416218 586442 416454
rect 586678 416218 586860 416454
rect 586260 416134 586860 416218
rect 586260 415898 586442 416134
rect 586678 415898 586860 416134
rect 586260 380454 586860 415898
rect 586260 380218 586442 380454
rect 586678 380218 586860 380454
rect 586260 380134 586860 380218
rect 586260 379898 586442 380134
rect 586678 379898 586860 380134
rect 586260 344454 586860 379898
rect 586260 344218 586442 344454
rect 586678 344218 586860 344454
rect 586260 344134 586860 344218
rect 586260 343898 586442 344134
rect 586678 343898 586860 344134
rect 586260 308454 586860 343898
rect 586260 308218 586442 308454
rect 586678 308218 586860 308454
rect 586260 308134 586860 308218
rect 586260 307898 586442 308134
rect 586678 307898 586860 308134
rect 586260 272454 586860 307898
rect 586260 272218 586442 272454
rect 586678 272218 586860 272454
rect 586260 272134 586860 272218
rect 586260 271898 586442 272134
rect 586678 271898 586860 272134
rect 586260 236454 586860 271898
rect 586260 236218 586442 236454
rect 586678 236218 586860 236454
rect 586260 236134 586860 236218
rect 586260 235898 586442 236134
rect 586678 235898 586860 236134
rect 586260 200454 586860 235898
rect 586260 200218 586442 200454
rect 586678 200218 586860 200454
rect 586260 200134 586860 200218
rect 586260 199898 586442 200134
rect 586678 199898 586860 200134
rect 586260 164454 586860 199898
rect 586260 164218 586442 164454
rect 586678 164218 586860 164454
rect 586260 164134 586860 164218
rect 586260 163898 586442 164134
rect 586678 163898 586860 164134
rect 586260 128454 586860 163898
rect 586260 128218 586442 128454
rect 586678 128218 586860 128454
rect 586260 128134 586860 128218
rect 586260 127898 586442 128134
rect 586678 127898 586860 128134
rect 586260 92454 586860 127898
rect 586260 92218 586442 92454
rect 586678 92218 586860 92454
rect 586260 92134 586860 92218
rect 586260 91898 586442 92134
rect 586678 91898 586860 92134
rect 586260 56454 586860 91898
rect 586260 56218 586442 56454
rect 586678 56218 586860 56454
rect 586260 56134 586860 56218
rect 586260 55898 586442 56134
rect 586678 55898 586860 56134
rect 586260 20454 586860 55898
rect 586260 20218 586442 20454
rect 586678 20218 586860 20454
rect 586260 20134 586860 20218
rect 586260 19898 586442 20134
rect 586678 19898 586860 20134
rect 586260 -1286 586860 19898
rect 586260 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect 586260 -1606 586860 -1522
rect 586260 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect 586260 -1864 586860 -1842
rect -3876 -2462 -3694 -2226
rect -3458 -2462 -3276 -2226
rect -3876 -2546 -3276 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 -3276 -2546
rect -3876 -2804 -3276 -2782
rect 587200 -2226 587800 706162
rect 587200 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect 587200 -2546 587800 -2462
rect 587200 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect 587200 -2804 587800 -2782
rect -4816 -3402 -4634 -3166
rect -4398 -3402 -4216 -3166
rect -4816 -3486 -4216 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 -4216 -3486
rect -4816 -3744 -4216 -3722
rect 588140 -3166 588740 707102
rect 588140 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect 588140 -3486 588740 -3402
rect 588140 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect 588140 -3744 588740 -3722
rect -5756 -4342 -5574 -4106
rect -5338 -4342 -5156 -4106
rect -5756 -4426 -5156 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 -5156 -4426
rect -5756 -4684 -5156 -4662
rect 589080 -4106 589680 708042
rect 589080 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect 589080 -4426 589680 -4342
rect 589080 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect 589080 -4684 589680 -4662
rect -6696 -5282 -6514 -5046
rect -6278 -5282 -6096 -5046
rect -6696 -5366 -6096 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 -6096 -5366
rect -6696 -5624 -6096 -5602
rect 590020 -5046 590620 708982
rect 590020 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect 590020 -5366 590620 -5282
rect 590020 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect 590020 -5624 590620 -5602
rect -7636 -6222 -7454 -5986
rect -7218 -6222 -7036 -5986
rect -7636 -6306 -7036 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 -7036 -6306
rect -7636 -6564 -7036 -6542
rect 590960 -5986 591560 709922
rect 590960 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect 590960 -6306 591560 -6222
rect 590960 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect 590960 -6564 591560 -6542
rect -8576 -7162 -8394 -6926
rect -8158 -7162 -7976 -6926
rect -8576 -7246 -7976 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 -7976 -7246
rect -8576 -7504 -7976 -7482
rect 591900 -6926 592500 710862
rect 591900 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect 591900 -7246 592500 -7162
rect 591900 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect 591900 -7504 592500 -7482
<< via4 >>
rect -8394 711182 -8158 711418
rect -8394 710862 -8158 711098
rect 592082 711182 592318 711418
rect 592082 710862 592318 711098
rect -7454 710242 -7218 710478
rect -7454 709922 -7218 710158
rect 591142 710242 591378 710478
rect 591142 709922 591378 710158
rect -6514 709302 -6278 709538
rect -6514 708982 -6278 709218
rect 590202 709302 590438 709538
rect 590202 708982 590438 709218
rect -5574 708362 -5338 708598
rect -5574 708042 -5338 708278
rect 589262 708362 589498 708598
rect 589262 708042 589498 708278
rect -4634 707422 -4398 707658
rect -4634 707102 -4398 707338
rect 588322 707422 588558 707658
rect 588322 707102 588558 707338
rect -3694 706482 -3458 706718
rect -3694 706162 -3458 706398
rect 587382 706482 587618 706718
rect 587382 706162 587618 706398
rect -2754 705542 -2518 705778
rect -2754 705222 -2518 705458
rect -2754 668218 -2518 668454
rect -2754 667898 -2518 668134
rect -2754 632218 -2518 632454
rect -2754 631898 -2518 632134
rect -2754 596218 -2518 596454
rect -2754 595898 -2518 596134
rect -2754 560218 -2518 560454
rect -2754 559898 -2518 560134
rect -2754 524218 -2518 524454
rect -2754 523898 -2518 524134
rect -2754 488218 -2518 488454
rect -2754 487898 -2518 488134
rect -2754 452218 -2518 452454
rect -2754 451898 -2518 452134
rect -2754 416218 -2518 416454
rect -2754 415898 -2518 416134
rect -2754 380218 -2518 380454
rect -2754 379898 -2518 380134
rect -2754 344218 -2518 344454
rect -2754 343898 -2518 344134
rect -2754 308218 -2518 308454
rect -2754 307898 -2518 308134
rect -2754 272218 -2518 272454
rect -2754 271898 -2518 272134
rect -2754 236218 -2518 236454
rect -2754 235898 -2518 236134
rect -2754 200218 -2518 200454
rect -2754 199898 -2518 200134
rect -2754 164218 -2518 164454
rect -2754 163898 -2518 164134
rect -2754 128218 -2518 128454
rect -2754 127898 -2518 128134
rect -2754 92218 -2518 92454
rect -2754 91898 -2518 92134
rect -2754 56218 -2518 56454
rect -2754 55898 -2518 56134
rect -2754 20218 -2518 20454
rect -2754 19898 -2518 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2754 -1522 -2518 -1286
rect -2754 -1842 -2518 -1606
rect 18986 705542 19222 705778
rect 18986 705222 19222 705458
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 54986 705542 55222 705778
rect 54986 705222 55222 705458
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 72986 614218 73222 614454
rect 72986 613898 73222 614134
rect 90986 705542 91222 705778
rect 90986 705222 91222 705458
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 90986 632218 91222 632454
rect 90986 631898 91222 632134
rect 90986 596218 91222 596454
rect 90986 595898 91222 596134
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 108986 614218 109222 614454
rect 108986 613898 109222 614134
rect 126986 705542 127222 705778
rect 126986 705222 127222 705458
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 126986 632218 127222 632454
rect 126986 631898 127222 632134
rect 126986 596218 127222 596454
rect 126986 595898 127222 596134
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 162986 705542 163222 705778
rect 162986 705222 163222 705458
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 198986 705542 199222 705778
rect 198986 705222 199222 705458
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 198986 632218 199222 632454
rect 198986 631898 199222 632134
rect 198986 596218 199222 596454
rect 198986 595898 199222 596134
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 216986 614218 217222 614454
rect 216986 613898 217222 614134
rect 234986 705542 235222 705778
rect 234986 705222 235222 705458
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 234986 632218 235222 632454
rect 234986 631898 235222 632134
rect 234986 596218 235222 596454
rect 234986 595898 235222 596134
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 252986 614218 253222 614454
rect 252986 613898 253222 614134
rect 270986 705542 271222 705778
rect 270986 705222 271222 705458
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 270986 596218 271222 596454
rect 270986 595898 271222 596134
rect 47130 578218 47366 578454
rect 47130 577898 47366 578134
rect 77850 578218 78086 578454
rect 77850 577898 78086 578134
rect 108570 578218 108806 578454
rect 108570 577898 108806 578134
rect 139290 578218 139526 578454
rect 139290 577898 139526 578134
rect 170010 578218 170246 578454
rect 170010 577898 170246 578134
rect 200730 578218 200966 578454
rect 200730 577898 200966 578134
rect 231450 578218 231686 578454
rect 231450 577898 231686 578134
rect 262170 578218 262406 578454
rect 262170 577898 262406 578134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 31770 560218 32006 560454
rect 31770 559898 32006 560134
rect 62490 560218 62726 560454
rect 62490 559898 62726 560134
rect 93210 560218 93446 560454
rect 93210 559898 93446 560134
rect 123930 560218 124166 560454
rect 123930 559898 124166 560134
rect 154650 560218 154886 560454
rect 154650 559898 154886 560134
rect 185370 560218 185606 560454
rect 185370 559898 185606 560134
rect 216090 560218 216326 560454
rect 216090 559898 216326 560134
rect 246810 560218 247046 560454
rect 246810 559898 247046 560134
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 47130 542218 47366 542454
rect 47130 541898 47366 542134
rect 77850 542218 78086 542454
rect 77850 541898 78086 542134
rect 108570 542218 108806 542454
rect 108570 541898 108806 542134
rect 139290 542218 139526 542454
rect 139290 541898 139526 542134
rect 170010 542218 170246 542454
rect 170010 541898 170246 542134
rect 200730 542218 200966 542454
rect 200730 541898 200966 542134
rect 231450 542218 231686 542454
rect 231450 541898 231686 542134
rect 262170 542218 262406 542454
rect 262170 541898 262406 542134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 31770 524218 32006 524454
rect 31770 523898 32006 524134
rect 62490 524218 62726 524454
rect 62490 523898 62726 524134
rect 93210 524218 93446 524454
rect 93210 523898 93446 524134
rect 123930 524218 124166 524454
rect 123930 523898 124166 524134
rect 154650 524218 154886 524454
rect 154650 523898 154886 524134
rect 185370 524218 185606 524454
rect 185370 523898 185606 524134
rect 216090 524218 216326 524454
rect 216090 523898 216326 524134
rect 246810 524218 247046 524454
rect 246810 523898 247046 524134
rect 270986 524218 271222 524454
rect 270986 523898 271222 524134
rect 47130 506218 47366 506454
rect 47130 505898 47366 506134
rect 77850 506218 78086 506454
rect 77850 505898 78086 506134
rect 108570 506218 108806 506454
rect 108570 505898 108806 506134
rect 139290 506218 139526 506454
rect 139290 505898 139526 506134
rect 170010 506218 170246 506454
rect 170010 505898 170246 506134
rect 200730 506218 200966 506454
rect 200730 505898 200966 506134
rect 231450 506218 231686 506454
rect 231450 505898 231686 506134
rect 262170 506218 262406 506454
rect 262170 505898 262406 506134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 31770 488218 32006 488454
rect 31770 487898 32006 488134
rect 62490 488218 62726 488454
rect 62490 487898 62726 488134
rect 93210 488218 93446 488454
rect 93210 487898 93446 488134
rect 123930 488218 124166 488454
rect 123930 487898 124166 488134
rect 154650 488218 154886 488454
rect 154650 487898 154886 488134
rect 185370 488218 185606 488454
rect 185370 487898 185606 488134
rect 216090 488218 216326 488454
rect 216090 487898 216326 488134
rect 246810 488218 247046 488454
rect 246810 487898 247046 488134
rect 270986 488218 271222 488454
rect 270986 487898 271222 488134
rect 47130 470218 47366 470454
rect 47130 469898 47366 470134
rect 77850 470218 78086 470454
rect 77850 469898 78086 470134
rect 108570 470218 108806 470454
rect 108570 469898 108806 470134
rect 139290 470218 139526 470454
rect 139290 469898 139526 470134
rect 170010 470218 170246 470454
rect 170010 469898 170246 470134
rect 200730 470218 200966 470454
rect 200730 469898 200966 470134
rect 231450 470218 231686 470454
rect 231450 469898 231686 470134
rect 262170 470218 262406 470454
rect 262170 469898 262406 470134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 31770 452218 32006 452454
rect 31770 451898 32006 452134
rect 62490 452218 62726 452454
rect 62490 451898 62726 452134
rect 93210 452218 93446 452454
rect 93210 451898 93446 452134
rect 123930 452218 124166 452454
rect 123930 451898 124166 452134
rect 154650 452218 154886 452454
rect 154650 451898 154886 452134
rect 185370 452218 185606 452454
rect 185370 451898 185606 452134
rect 216090 452218 216326 452454
rect 216090 451898 216326 452134
rect 246810 452218 247046 452454
rect 246810 451898 247046 452134
rect 270986 452218 271222 452454
rect 270986 451898 271222 452134
rect 47130 434218 47366 434454
rect 47130 433898 47366 434134
rect 77850 434218 78086 434454
rect 77850 433898 78086 434134
rect 108570 434218 108806 434454
rect 108570 433898 108806 434134
rect 139290 434218 139526 434454
rect 139290 433898 139526 434134
rect 170010 434218 170246 434454
rect 170010 433898 170246 434134
rect 200730 434218 200966 434454
rect 200730 433898 200966 434134
rect 231450 434218 231686 434454
rect 231450 433898 231686 434134
rect 262170 434218 262406 434454
rect 262170 433898 262406 434134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 31770 416218 32006 416454
rect 31770 415898 32006 416134
rect 62490 416218 62726 416454
rect 62490 415898 62726 416134
rect 93210 416218 93446 416454
rect 93210 415898 93446 416134
rect 123930 416218 124166 416454
rect 123930 415898 124166 416134
rect 154650 416218 154886 416454
rect 154650 415898 154886 416134
rect 185370 416218 185606 416454
rect 185370 415898 185606 416134
rect 216090 416218 216326 416454
rect 216090 415898 216326 416134
rect 246810 416218 247046 416454
rect 246810 415898 247046 416134
rect 270986 416218 271222 416454
rect 270986 415898 271222 416134
rect 47130 398218 47366 398454
rect 47130 397898 47366 398134
rect 77850 398218 78086 398454
rect 77850 397898 78086 398134
rect 108570 398218 108806 398454
rect 108570 397898 108806 398134
rect 139290 398218 139526 398454
rect 139290 397898 139526 398134
rect 170010 398218 170246 398454
rect 170010 397898 170246 398134
rect 200730 398218 200966 398454
rect 200730 397898 200966 398134
rect 231450 398218 231686 398454
rect 231450 397898 231686 398134
rect 262170 398218 262406 398454
rect 262170 397898 262406 398134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 72986 362218 73222 362454
rect 72986 361898 73222 362134
rect 72986 326218 73222 326454
rect 72986 325898 73222 326134
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 90986 380218 91222 380454
rect 90986 379898 91222 380134
rect 90986 344218 91222 344454
rect 90986 343898 91222 344134
rect 90986 308218 91222 308454
rect 90986 307898 91222 308134
rect 108986 362218 109222 362454
rect 108986 361898 109222 362134
rect 108986 326218 109222 326454
rect 108986 325898 109222 326134
rect 108986 290218 109222 290454
rect 108986 289898 109222 290134
rect 126986 380218 127222 380454
rect 126986 379898 127222 380134
rect 126986 344218 127222 344454
rect 126986 343898 127222 344134
rect 126986 308218 127222 308454
rect 126986 307898 127222 308134
rect 144986 362218 145222 362454
rect 144986 361898 145222 362134
rect 144986 326218 145222 326454
rect 144986 325898 145222 326134
rect 144986 290218 145222 290454
rect 144986 289898 145222 290134
rect 162986 380218 163222 380454
rect 162986 379898 163222 380134
rect 162986 344218 163222 344454
rect 162986 343898 163222 344134
rect 162986 308218 163222 308454
rect 162986 307898 163222 308134
rect 180986 362218 181222 362454
rect 180986 361898 181222 362134
rect 180986 326218 181222 326454
rect 180986 325898 181222 326134
rect 180986 290218 181222 290454
rect 180986 289898 181222 290134
rect 198986 380218 199222 380454
rect 198986 379898 199222 380134
rect 198986 344218 199222 344454
rect 198986 343898 199222 344134
rect 198986 308218 199222 308454
rect 198986 307898 199222 308134
rect 216986 362218 217222 362454
rect 216986 361898 217222 362134
rect 216986 326218 217222 326454
rect 216986 325898 217222 326134
rect 216986 290218 217222 290454
rect 216986 289898 217222 290134
rect 234986 380218 235222 380454
rect 234986 379898 235222 380134
rect 234986 344218 235222 344454
rect 234986 343898 235222 344134
rect 234986 308218 235222 308454
rect 234986 307898 235222 308134
rect 252986 362218 253222 362454
rect 252986 361898 253222 362134
rect 270986 380218 271222 380454
rect 270986 379898 271222 380134
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 288986 542218 289222 542454
rect 288986 541898 289222 542134
rect 288986 506218 289222 506454
rect 288986 505898 289222 506134
rect 288986 470218 289222 470454
rect 288986 469898 289222 470134
rect 288986 434218 289222 434454
rect 288986 433898 289222 434134
rect 288986 398218 289222 398454
rect 288986 397898 289222 398134
rect 288986 362218 289222 362454
rect 288986 361898 289222 362134
rect 306986 705542 307222 705778
rect 306986 705222 307222 705458
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 306986 596218 307222 596454
rect 306986 595898 307222 596134
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 324986 650218 325222 650454
rect 324986 649898 325222 650134
rect 324986 614218 325222 614454
rect 324986 613898 325222 614134
rect 342986 705542 343222 705778
rect 342986 705222 343222 705458
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 342986 632218 343222 632454
rect 342986 631898 343222 632134
rect 342986 596218 343222 596454
rect 342986 595898 343222 596134
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 360986 650218 361222 650454
rect 360986 649898 361222 650134
rect 360986 614218 361222 614454
rect 360986 613898 361222 614134
rect 378986 705542 379222 705778
rect 378986 705222 379222 705458
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 378986 632218 379222 632454
rect 378986 631898 379222 632134
rect 378986 596218 379222 596454
rect 378986 595898 379222 596134
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 414986 705542 415222 705778
rect 414986 705222 415222 705458
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 414986 596218 415222 596454
rect 414986 595898 415222 596134
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 450986 705542 451222 705778
rect 450986 705222 451222 705458
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 450986 632218 451222 632454
rect 450986 631898 451222 632134
rect 450986 596218 451222 596454
rect 450986 595898 451222 596134
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 468986 614218 469222 614454
rect 468986 613898 469222 614134
rect 486986 705542 487222 705778
rect 486986 705222 487222 705458
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 486986 632218 487222 632454
rect 486986 631898 487222 632134
rect 486986 596218 487222 596454
rect 486986 595898 487222 596134
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 504986 614218 505222 614454
rect 504986 613898 505222 614134
rect 522986 705542 523222 705778
rect 522986 705222 523222 705458
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 558986 705542 559222 705778
rect 558986 705222 559222 705458
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 586442 705542 586678 705778
rect 586442 705222 586678 705458
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 339258 578218 339494 578454
rect 339258 577898 339494 578134
rect 369978 578218 370214 578454
rect 369978 577898 370214 578134
rect 400698 578218 400934 578454
rect 400698 577898 400934 578134
rect 431418 578218 431654 578454
rect 431418 577898 431654 578134
rect 462138 578218 462374 578454
rect 462138 577898 462374 578134
rect 492858 578218 493094 578454
rect 492858 577898 493094 578134
rect 523578 578218 523814 578454
rect 523578 577898 523814 578134
rect 554298 578218 554534 578454
rect 554298 577898 554534 578134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 306986 560218 307222 560454
rect 306986 559898 307222 560134
rect 323898 560218 324134 560454
rect 323898 559898 324134 560134
rect 354618 560218 354854 560454
rect 354618 559898 354854 560134
rect 385338 560218 385574 560454
rect 385338 559898 385574 560134
rect 416058 560218 416294 560454
rect 416058 559898 416294 560134
rect 446778 560218 447014 560454
rect 446778 559898 447014 560134
rect 477498 560218 477734 560454
rect 477498 559898 477734 560134
rect 508218 560218 508454 560454
rect 508218 559898 508454 560134
rect 538938 560218 539174 560454
rect 538938 559898 539174 560134
rect 339258 542218 339494 542454
rect 339258 541898 339494 542134
rect 369978 542218 370214 542454
rect 369978 541898 370214 542134
rect 400698 542218 400934 542454
rect 400698 541898 400934 542134
rect 431418 542218 431654 542454
rect 431418 541898 431654 542134
rect 462138 542218 462374 542454
rect 462138 541898 462374 542134
rect 492858 542218 493094 542454
rect 492858 541898 493094 542134
rect 523578 542218 523814 542454
rect 523578 541898 523814 542134
rect 554298 542218 554534 542454
rect 554298 541898 554534 542134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 306986 524218 307222 524454
rect 306986 523898 307222 524134
rect 323898 524218 324134 524454
rect 323898 523898 324134 524134
rect 354618 524218 354854 524454
rect 354618 523898 354854 524134
rect 385338 524218 385574 524454
rect 385338 523898 385574 524134
rect 416058 524218 416294 524454
rect 416058 523898 416294 524134
rect 446778 524218 447014 524454
rect 446778 523898 447014 524134
rect 477498 524218 477734 524454
rect 477498 523898 477734 524134
rect 508218 524218 508454 524454
rect 508218 523898 508454 524134
rect 538938 524218 539174 524454
rect 538938 523898 539174 524134
rect 339258 506218 339494 506454
rect 339258 505898 339494 506134
rect 369978 506218 370214 506454
rect 369978 505898 370214 506134
rect 400698 506218 400934 506454
rect 400698 505898 400934 506134
rect 431418 506218 431654 506454
rect 431418 505898 431654 506134
rect 462138 506218 462374 506454
rect 462138 505898 462374 506134
rect 492858 506218 493094 506454
rect 492858 505898 493094 506134
rect 523578 506218 523814 506454
rect 523578 505898 523814 506134
rect 554298 506218 554534 506454
rect 554298 505898 554534 506134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 306986 488218 307222 488454
rect 306986 487898 307222 488134
rect 323898 488218 324134 488454
rect 323898 487898 324134 488134
rect 354618 488218 354854 488454
rect 354618 487898 354854 488134
rect 385338 488218 385574 488454
rect 385338 487898 385574 488134
rect 416058 488218 416294 488454
rect 416058 487898 416294 488134
rect 446778 488218 447014 488454
rect 446778 487898 447014 488134
rect 477498 488218 477734 488454
rect 477498 487898 477734 488134
rect 508218 488218 508454 488454
rect 508218 487898 508454 488134
rect 538938 488218 539174 488454
rect 538938 487898 539174 488134
rect 339258 470218 339494 470454
rect 339258 469898 339494 470134
rect 369978 470218 370214 470454
rect 369978 469898 370214 470134
rect 400698 470218 400934 470454
rect 400698 469898 400934 470134
rect 431418 470218 431654 470454
rect 431418 469898 431654 470134
rect 462138 470218 462374 470454
rect 462138 469898 462374 470134
rect 492858 470218 493094 470454
rect 492858 469898 493094 470134
rect 523578 470218 523814 470454
rect 523578 469898 523814 470134
rect 554298 470218 554534 470454
rect 554298 469898 554534 470134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 306986 452218 307222 452454
rect 306986 451898 307222 452134
rect 323898 452218 324134 452454
rect 323898 451898 324134 452134
rect 354618 452218 354854 452454
rect 354618 451898 354854 452134
rect 385338 452218 385574 452454
rect 385338 451898 385574 452134
rect 416058 452218 416294 452454
rect 416058 451898 416294 452134
rect 446778 452218 447014 452454
rect 446778 451898 447014 452134
rect 477498 452218 477734 452454
rect 477498 451898 477734 452134
rect 508218 452218 508454 452454
rect 508218 451898 508454 452134
rect 538938 452218 539174 452454
rect 538938 451898 539174 452134
rect 339258 434218 339494 434454
rect 339258 433898 339494 434134
rect 369978 434218 370214 434454
rect 369978 433898 370214 434134
rect 400698 434218 400934 434454
rect 400698 433898 400934 434134
rect 431418 434218 431654 434454
rect 431418 433898 431654 434134
rect 462138 434218 462374 434454
rect 462138 433898 462374 434134
rect 492858 434218 493094 434454
rect 492858 433898 493094 434134
rect 523578 434218 523814 434454
rect 523578 433898 523814 434134
rect 554298 434218 554534 434454
rect 554298 433898 554534 434134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 306986 416218 307222 416454
rect 306986 415898 307222 416134
rect 323898 416218 324134 416454
rect 323898 415898 324134 416134
rect 354618 416218 354854 416454
rect 354618 415898 354854 416134
rect 385338 416218 385574 416454
rect 385338 415898 385574 416134
rect 416058 416218 416294 416454
rect 416058 415898 416294 416134
rect 446778 416218 447014 416454
rect 446778 415898 447014 416134
rect 477498 416218 477734 416454
rect 477498 415898 477734 416134
rect 508218 416218 508454 416454
rect 508218 415898 508454 416134
rect 538938 416218 539174 416454
rect 538938 415898 539174 416134
rect 339258 398218 339494 398454
rect 339258 397898 339494 398134
rect 369978 398218 370214 398454
rect 369978 397898 370214 398134
rect 400698 398218 400934 398454
rect 400698 397898 400934 398134
rect 431418 398218 431654 398454
rect 431418 397898 431654 398134
rect 462138 398218 462374 398454
rect 462138 397898 462374 398134
rect 492858 398218 493094 398454
rect 492858 397898 493094 398134
rect 523578 398218 523814 398454
rect 523578 397898 523814 398134
rect 554298 398218 554534 398454
rect 554298 397898 554534 398134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 306986 380218 307222 380454
rect 306986 379898 307222 380134
rect 324986 362218 325222 362454
rect 324986 361898 325222 362134
rect 292154 344218 292390 344454
rect 292154 343898 292390 344134
rect 252986 326218 253222 326454
rect 252986 325898 253222 326134
rect 276794 326218 277030 326454
rect 276794 325898 277030 326134
rect 307514 326218 307750 326454
rect 307514 325898 307750 326134
rect 324986 326218 325222 326454
rect 324986 325898 325222 326134
rect 252986 290218 253222 290454
rect 252986 289898 253222 290134
rect 270986 308218 271222 308454
rect 270986 307898 271222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 270986 272218 271222 272454
rect 270986 271898 271222 272134
rect 47130 254218 47366 254454
rect 47130 253898 47366 254134
rect 77850 254218 78086 254454
rect 77850 253898 78086 254134
rect 108570 254218 108806 254454
rect 108570 253898 108806 254134
rect 139290 254218 139526 254454
rect 139290 253898 139526 254134
rect 170010 254218 170246 254454
rect 170010 253898 170246 254134
rect 200730 254218 200966 254454
rect 200730 253898 200966 254134
rect 231450 254218 231686 254454
rect 231450 253898 231686 254134
rect 262170 254218 262406 254454
rect 262170 253898 262406 254134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 31770 236218 32006 236454
rect 31770 235898 32006 236134
rect 62490 236218 62726 236454
rect 62490 235898 62726 236134
rect 93210 236218 93446 236454
rect 93210 235898 93446 236134
rect 123930 236218 124166 236454
rect 123930 235898 124166 236134
rect 154650 236218 154886 236454
rect 154650 235898 154886 236134
rect 185370 236218 185606 236454
rect 185370 235898 185606 236134
rect 216090 236218 216326 236454
rect 216090 235898 216326 236134
rect 246810 236218 247046 236454
rect 246810 235898 247046 236134
rect 270986 236218 271222 236454
rect 270986 235898 271222 236134
rect 47130 218218 47366 218454
rect 47130 217898 47366 218134
rect 77850 218218 78086 218454
rect 77850 217898 78086 218134
rect 108570 218218 108806 218454
rect 108570 217898 108806 218134
rect 139290 218218 139526 218454
rect 139290 217898 139526 218134
rect 170010 218218 170246 218454
rect 170010 217898 170246 218134
rect 200730 218218 200966 218454
rect 200730 217898 200966 218134
rect 231450 218218 231686 218454
rect 231450 217898 231686 218134
rect 262170 218218 262406 218454
rect 262170 217898 262406 218134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 31770 200218 32006 200454
rect 31770 199898 32006 200134
rect 62490 200218 62726 200454
rect 62490 199898 62726 200134
rect 93210 200218 93446 200454
rect 93210 199898 93446 200134
rect 123930 200218 124166 200454
rect 123930 199898 124166 200134
rect 154650 200218 154886 200454
rect 154650 199898 154886 200134
rect 185370 200218 185606 200454
rect 185370 199898 185606 200134
rect 216090 200218 216326 200454
rect 216090 199898 216326 200134
rect 246810 200218 247046 200454
rect 246810 199898 247046 200134
rect 270986 200218 271222 200454
rect 270986 199898 271222 200134
rect 47130 182218 47366 182454
rect 47130 181898 47366 182134
rect 77850 182218 78086 182454
rect 77850 181898 78086 182134
rect 108570 182218 108806 182454
rect 108570 181898 108806 182134
rect 139290 182218 139526 182454
rect 139290 181898 139526 182134
rect 170010 182218 170246 182454
rect 170010 181898 170246 182134
rect 200730 182218 200966 182454
rect 200730 181898 200966 182134
rect 231450 182218 231686 182454
rect 231450 181898 231686 182134
rect 262170 182218 262406 182454
rect 262170 181898 262406 182134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 31770 164218 32006 164454
rect 31770 163898 32006 164134
rect 62490 164218 62726 164454
rect 62490 163898 62726 164134
rect 93210 164218 93446 164454
rect 93210 163898 93446 164134
rect 123930 164218 124166 164454
rect 123930 163898 124166 164134
rect 154650 164218 154886 164454
rect 154650 163898 154886 164134
rect 185370 164218 185606 164454
rect 185370 163898 185606 164134
rect 216090 164218 216326 164454
rect 216090 163898 216326 164134
rect 246810 164218 247046 164454
rect 246810 163898 247046 164134
rect 270986 164218 271222 164454
rect 270986 163898 271222 164134
rect 47130 146218 47366 146454
rect 47130 145898 47366 146134
rect 77850 146218 78086 146454
rect 77850 145898 78086 146134
rect 108570 146218 108806 146454
rect 108570 145898 108806 146134
rect 139290 146218 139526 146454
rect 139290 145898 139526 146134
rect 170010 146218 170246 146454
rect 170010 145898 170246 146134
rect 200730 146218 200966 146454
rect 200730 145898 200966 146134
rect 231450 146218 231686 146454
rect 231450 145898 231686 146134
rect 262170 146218 262406 146454
rect 262170 145898 262406 146134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 31770 128218 32006 128454
rect 31770 127898 32006 128134
rect 62490 128218 62726 128454
rect 62490 127898 62726 128134
rect 93210 128218 93446 128454
rect 93210 127898 93446 128134
rect 123930 128218 124166 128454
rect 123930 127898 124166 128134
rect 154650 128218 154886 128454
rect 154650 127898 154886 128134
rect 185370 128218 185606 128454
rect 185370 127898 185606 128134
rect 216090 128218 216326 128454
rect 216090 127898 216326 128134
rect 246810 128218 247046 128454
rect 246810 127898 247046 128134
rect 270986 128218 271222 128454
rect 270986 127898 271222 128134
rect 47130 110218 47366 110454
rect 47130 109898 47366 110134
rect 77850 110218 78086 110454
rect 77850 109898 78086 110134
rect 108570 110218 108806 110454
rect 108570 109898 108806 110134
rect 139290 110218 139526 110454
rect 139290 109898 139526 110134
rect 170010 110218 170246 110454
rect 170010 109898 170246 110134
rect 200730 110218 200966 110454
rect 200730 109898 200966 110134
rect 231450 110218 231686 110454
rect 231450 109898 231686 110134
rect 262170 110218 262406 110454
rect 262170 109898 262406 110134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 31770 92218 32006 92454
rect 31770 91898 32006 92134
rect 62490 92218 62726 92454
rect 62490 91898 62726 92134
rect 93210 92218 93446 92454
rect 93210 91898 93446 92134
rect 123930 92218 124166 92454
rect 123930 91898 124166 92134
rect 154650 92218 154886 92454
rect 154650 91898 154886 92134
rect 185370 92218 185606 92454
rect 185370 91898 185606 92134
rect 216090 92218 216326 92454
rect 216090 91898 216326 92134
rect 246810 92218 247046 92454
rect 246810 91898 247046 92134
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1522 19222 -1286
rect 18986 -1842 19222 -1606
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1522 55222 -1286
rect 54986 -1842 55222 -1606
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1522 91222 -1286
rect 90986 -1842 91222 -1606
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1522 127222 -1286
rect 126986 -1842 127222 -1606
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1522 163222 -1286
rect 162986 -1842 163222 -1606
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1522 199222 -1286
rect 198986 -1842 199222 -1606
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1522 235222 -1286
rect 234986 -1842 235222 -1606
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1522 271222 -1286
rect 270986 -1842 271222 -1606
rect 288986 290218 289222 290454
rect 288986 289898 289222 290134
rect 288986 254218 289222 254454
rect 288986 253898 289222 254134
rect 288986 218218 289222 218454
rect 288986 217898 289222 218134
rect 288986 182218 289222 182454
rect 288986 181898 289222 182134
rect 288986 146218 289222 146454
rect 288986 145898 289222 146134
rect 288986 110218 289222 110454
rect 288986 109898 289222 110134
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 306986 308218 307222 308454
rect 306986 307898 307222 308134
rect 324986 290218 325222 290454
rect 324986 289898 325222 290134
rect 342986 380218 343222 380454
rect 342986 379898 343222 380134
rect 342986 344218 343222 344454
rect 342986 343898 343222 344134
rect 342986 308218 343222 308454
rect 342986 307898 343222 308134
rect 360986 362218 361222 362454
rect 360986 361898 361222 362134
rect 360986 326218 361222 326454
rect 360986 325898 361222 326134
rect 360986 290218 361222 290454
rect 360986 289898 361222 290134
rect 378986 380218 379222 380454
rect 378986 379898 379222 380134
rect 378986 344218 379222 344454
rect 378986 343898 379222 344134
rect 378986 308218 379222 308454
rect 378986 307898 379222 308134
rect 396986 362218 397222 362454
rect 396986 361898 397222 362134
rect 396986 326218 397222 326454
rect 396986 325898 397222 326134
rect 396986 290218 397222 290454
rect 396986 289898 397222 290134
rect 414986 380218 415222 380454
rect 414986 379898 415222 380134
rect 414986 344218 415222 344454
rect 414986 343898 415222 344134
rect 414986 308218 415222 308454
rect 414986 307898 415222 308134
rect 432986 362218 433222 362454
rect 432986 361898 433222 362134
rect 432986 326218 433222 326454
rect 432986 325898 433222 326134
rect 432986 290218 433222 290454
rect 432986 289898 433222 290134
rect 450986 380218 451222 380454
rect 450986 379898 451222 380134
rect 450986 344218 451222 344454
rect 450986 343898 451222 344134
rect 450986 308218 451222 308454
rect 450986 307898 451222 308134
rect 468986 362218 469222 362454
rect 468986 361898 469222 362134
rect 468986 326218 469222 326454
rect 468986 325898 469222 326134
rect 468986 290218 469222 290454
rect 468986 289898 469222 290134
rect 486986 380218 487222 380454
rect 486986 379898 487222 380134
rect 486986 344218 487222 344454
rect 486986 343898 487222 344134
rect 486986 308218 487222 308454
rect 486986 307898 487222 308134
rect 504986 362218 505222 362454
rect 504986 361898 505222 362134
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 306986 272218 307222 272454
rect 306986 271898 307222 272134
rect 339258 254218 339494 254454
rect 339258 253898 339494 254134
rect 369978 254218 370214 254454
rect 369978 253898 370214 254134
rect 400698 254218 400934 254454
rect 400698 253898 400934 254134
rect 431418 254218 431654 254454
rect 431418 253898 431654 254134
rect 462138 254218 462374 254454
rect 462138 253898 462374 254134
rect 492858 254218 493094 254454
rect 492858 253898 493094 254134
rect 523578 254218 523814 254454
rect 523578 253898 523814 254134
rect 554298 254218 554534 254454
rect 554298 253898 554534 254134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 306986 236218 307222 236454
rect 306986 235898 307222 236134
rect 323898 236218 324134 236454
rect 323898 235898 324134 236134
rect 354618 236218 354854 236454
rect 354618 235898 354854 236134
rect 385338 236218 385574 236454
rect 385338 235898 385574 236134
rect 416058 236218 416294 236454
rect 416058 235898 416294 236134
rect 446778 236218 447014 236454
rect 446778 235898 447014 236134
rect 477498 236218 477734 236454
rect 477498 235898 477734 236134
rect 508218 236218 508454 236454
rect 508218 235898 508454 236134
rect 538938 236218 539174 236454
rect 538938 235898 539174 236134
rect 339258 218218 339494 218454
rect 339258 217898 339494 218134
rect 369978 218218 370214 218454
rect 369978 217898 370214 218134
rect 400698 218218 400934 218454
rect 400698 217898 400934 218134
rect 431418 218218 431654 218454
rect 431418 217898 431654 218134
rect 462138 218218 462374 218454
rect 462138 217898 462374 218134
rect 492858 218218 493094 218454
rect 492858 217898 493094 218134
rect 523578 218218 523814 218454
rect 523578 217898 523814 218134
rect 554298 218218 554534 218454
rect 554298 217898 554534 218134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 306986 200218 307222 200454
rect 306986 199898 307222 200134
rect 323898 200218 324134 200454
rect 323898 199898 324134 200134
rect 354618 200218 354854 200454
rect 354618 199898 354854 200134
rect 385338 200218 385574 200454
rect 385338 199898 385574 200134
rect 416058 200218 416294 200454
rect 416058 199898 416294 200134
rect 446778 200218 447014 200454
rect 446778 199898 447014 200134
rect 477498 200218 477734 200454
rect 477498 199898 477734 200134
rect 508218 200218 508454 200454
rect 508218 199898 508454 200134
rect 538938 200218 539174 200454
rect 538938 199898 539174 200134
rect 339258 182218 339494 182454
rect 339258 181898 339494 182134
rect 369978 182218 370214 182454
rect 369978 181898 370214 182134
rect 400698 182218 400934 182454
rect 400698 181898 400934 182134
rect 431418 182218 431654 182454
rect 431418 181898 431654 182134
rect 462138 182218 462374 182454
rect 462138 181898 462374 182134
rect 492858 182218 493094 182454
rect 492858 181898 493094 182134
rect 523578 182218 523814 182454
rect 523578 181898 523814 182134
rect 554298 182218 554534 182454
rect 554298 181898 554534 182134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 306986 164218 307222 164454
rect 306986 163898 307222 164134
rect 323898 164218 324134 164454
rect 323898 163898 324134 164134
rect 354618 164218 354854 164454
rect 354618 163898 354854 164134
rect 385338 164218 385574 164454
rect 385338 163898 385574 164134
rect 416058 164218 416294 164454
rect 416058 163898 416294 164134
rect 446778 164218 447014 164454
rect 446778 163898 447014 164134
rect 477498 164218 477734 164454
rect 477498 163898 477734 164134
rect 508218 164218 508454 164454
rect 508218 163898 508454 164134
rect 538938 164218 539174 164454
rect 538938 163898 539174 164134
rect 339258 146218 339494 146454
rect 339258 145898 339494 146134
rect 369978 146218 370214 146454
rect 369978 145898 370214 146134
rect 400698 146218 400934 146454
rect 400698 145898 400934 146134
rect 431418 146218 431654 146454
rect 431418 145898 431654 146134
rect 462138 146218 462374 146454
rect 462138 145898 462374 146134
rect 492858 146218 493094 146454
rect 492858 145898 493094 146134
rect 523578 146218 523814 146454
rect 523578 145898 523814 146134
rect 554298 146218 554534 146454
rect 554298 145898 554534 146134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 306986 128218 307222 128454
rect 306986 127898 307222 128134
rect 323898 128218 324134 128454
rect 323898 127898 324134 128134
rect 354618 128218 354854 128454
rect 354618 127898 354854 128134
rect 385338 128218 385574 128454
rect 385338 127898 385574 128134
rect 416058 128218 416294 128454
rect 416058 127898 416294 128134
rect 446778 128218 447014 128454
rect 446778 127898 447014 128134
rect 477498 128218 477734 128454
rect 477498 127898 477734 128134
rect 508218 128218 508454 128454
rect 508218 127898 508454 128134
rect 538938 128218 539174 128454
rect 538938 127898 539174 128134
rect 339258 110218 339494 110454
rect 339258 109898 339494 110134
rect 369978 110218 370214 110454
rect 369978 109898 370214 110134
rect 400698 110218 400934 110454
rect 400698 109898 400934 110134
rect 431418 110218 431654 110454
rect 431418 109898 431654 110134
rect 462138 110218 462374 110454
rect 462138 109898 462374 110134
rect 492858 110218 493094 110454
rect 492858 109898 493094 110134
rect 523578 110218 523814 110454
rect 523578 109898 523814 110134
rect 554298 110218 554534 110454
rect 554298 109898 554534 110134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 323898 92218 324134 92454
rect 323898 91898 324134 92134
rect 354618 92218 354854 92454
rect 354618 91898 354854 92134
rect 385338 92218 385574 92454
rect 385338 91898 385574 92134
rect 416058 92218 416294 92454
rect 416058 91898 416294 92134
rect 446778 92218 447014 92454
rect 446778 91898 447014 92134
rect 477498 92218 477734 92454
rect 477498 91898 477734 92134
rect 508218 92218 508454 92454
rect 508218 91898 508454 92134
rect 538938 92218 539174 92454
rect 538938 91898 539174 92134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1522 307222 -1286
rect 306986 -1842 307222 -1606
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1522 343222 -1286
rect 342986 -1842 343222 -1606
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1522 379222 -1286
rect 378986 -1842 379222 -1606
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1522 415222 -1286
rect 414986 -1842 415222 -1606
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1522 451222 -1286
rect 450986 -1842 451222 -1606
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1522 487222 -1286
rect 486986 -1842 487222 -1606
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1522 523222 -1286
rect 522986 -1842 523222 -1606
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1522 559222 -1286
rect 558986 -1842 559222 -1606
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586442 668218 586678 668454
rect 586442 667898 586678 668134
rect 586442 632218 586678 632454
rect 586442 631898 586678 632134
rect 586442 596218 586678 596454
rect 586442 595898 586678 596134
rect 586442 560218 586678 560454
rect 586442 559898 586678 560134
rect 586442 524218 586678 524454
rect 586442 523898 586678 524134
rect 586442 488218 586678 488454
rect 586442 487898 586678 488134
rect 586442 452218 586678 452454
rect 586442 451898 586678 452134
rect 586442 416218 586678 416454
rect 586442 415898 586678 416134
rect 586442 380218 586678 380454
rect 586442 379898 586678 380134
rect 586442 344218 586678 344454
rect 586442 343898 586678 344134
rect 586442 308218 586678 308454
rect 586442 307898 586678 308134
rect 586442 272218 586678 272454
rect 586442 271898 586678 272134
rect 586442 236218 586678 236454
rect 586442 235898 586678 236134
rect 586442 200218 586678 200454
rect 586442 199898 586678 200134
rect 586442 164218 586678 164454
rect 586442 163898 586678 164134
rect 586442 128218 586678 128454
rect 586442 127898 586678 128134
rect 586442 92218 586678 92454
rect 586442 91898 586678 92134
rect 586442 56218 586678 56454
rect 586442 55898 586678 56134
rect 586442 20218 586678 20454
rect 586442 19898 586678 20134
rect 586442 -1522 586678 -1286
rect 586442 -1842 586678 -1606
rect -3694 -2462 -3458 -2226
rect -3694 -2782 -3458 -2546
rect 587382 -2462 587618 -2226
rect 587382 -2782 587618 -2546
rect -4634 -3402 -4398 -3166
rect -4634 -3722 -4398 -3486
rect 588322 -3402 588558 -3166
rect 588322 -3722 588558 -3486
rect -5574 -4342 -5338 -4106
rect -5574 -4662 -5338 -4426
rect 589262 -4342 589498 -4106
rect 589262 -4662 589498 -4426
rect -6514 -5282 -6278 -5046
rect -6514 -5602 -6278 -5366
rect 590202 -5282 590438 -5046
rect 590202 -5602 590438 -5366
rect -7454 -6222 -7218 -5986
rect -7454 -6542 -7218 -6306
rect 591142 -6222 591378 -5986
rect 591142 -6542 591378 -6306
rect -8394 -7162 -8158 -6926
rect -8394 -7482 -8158 -7246
rect 592082 -7162 592318 -6926
rect 592082 -7482 592318 -7246
<< metal5 >>
rect -8576 711440 -7976 711442
rect 591900 711440 592500 711442
rect -8576 711418 592500 711440
rect -8576 711182 -8394 711418
rect -8158 711182 592082 711418
rect 592318 711182 592500 711418
rect -8576 711098 592500 711182
rect -8576 710862 -8394 711098
rect -8158 710862 592082 711098
rect 592318 710862 592500 711098
rect -8576 710840 592500 710862
rect -8576 710838 -7976 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 590960 710500 591560 710502
rect -7636 710478 591560 710500
rect -7636 710242 -7454 710478
rect -7218 710242 591142 710478
rect 591378 710242 591560 710478
rect -7636 710158 591560 710242
rect -7636 709922 -7454 710158
rect -7218 709922 591142 710158
rect 591378 709922 591560 710158
rect -7636 709900 591560 709922
rect -7636 709898 -7036 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 590020 709560 590620 709562
rect -6696 709538 590620 709560
rect -6696 709302 -6514 709538
rect -6278 709302 590202 709538
rect 590438 709302 590620 709538
rect -6696 709218 590620 709302
rect -6696 708982 -6514 709218
rect -6278 708982 590202 709218
rect 590438 708982 590620 709218
rect -6696 708960 590620 708982
rect -6696 708958 -6096 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 589080 708620 589680 708622
rect -5756 708598 589680 708620
rect -5756 708362 -5574 708598
rect -5338 708362 589262 708598
rect 589498 708362 589680 708598
rect -5756 708278 589680 708362
rect -5756 708042 -5574 708278
rect -5338 708042 589262 708278
rect 589498 708042 589680 708278
rect -5756 708020 589680 708042
rect -5756 708018 -5156 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 588140 707680 588740 707682
rect -4816 707658 588740 707680
rect -4816 707422 -4634 707658
rect -4398 707422 588322 707658
rect 588558 707422 588740 707658
rect -4816 707338 588740 707422
rect -4816 707102 -4634 707338
rect -4398 707102 588322 707338
rect 588558 707102 588740 707338
rect -4816 707080 588740 707102
rect -4816 707078 -4216 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 587200 706740 587800 706742
rect -3876 706718 587800 706740
rect -3876 706482 -3694 706718
rect -3458 706482 587382 706718
rect 587618 706482 587800 706718
rect -3876 706398 587800 706482
rect -3876 706162 -3694 706398
rect -3458 706162 587382 706398
rect 587618 706162 587800 706398
rect -3876 706140 587800 706162
rect -3876 706138 -3276 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 18804 705800 19404 705802
rect 54804 705800 55404 705802
rect 90804 705800 91404 705802
rect 126804 705800 127404 705802
rect 162804 705800 163404 705802
rect 198804 705800 199404 705802
rect 234804 705800 235404 705802
rect 270804 705800 271404 705802
rect 306804 705800 307404 705802
rect 342804 705800 343404 705802
rect 378804 705800 379404 705802
rect 414804 705800 415404 705802
rect 450804 705800 451404 705802
rect 486804 705800 487404 705802
rect 522804 705800 523404 705802
rect 558804 705800 559404 705802
rect 586260 705800 586860 705802
rect -2936 705778 586860 705800
rect -2936 705542 -2754 705778
rect -2518 705542 18986 705778
rect 19222 705542 54986 705778
rect 55222 705542 90986 705778
rect 91222 705542 126986 705778
rect 127222 705542 162986 705778
rect 163222 705542 198986 705778
rect 199222 705542 234986 705778
rect 235222 705542 270986 705778
rect 271222 705542 306986 705778
rect 307222 705542 342986 705778
rect 343222 705542 378986 705778
rect 379222 705542 414986 705778
rect 415222 705542 450986 705778
rect 451222 705542 486986 705778
rect 487222 705542 522986 705778
rect 523222 705542 558986 705778
rect 559222 705542 586442 705778
rect 586678 705542 586860 705778
rect -2936 705458 586860 705542
rect -2936 705222 -2754 705458
rect -2518 705222 18986 705458
rect 19222 705222 54986 705458
rect 55222 705222 90986 705458
rect 91222 705222 126986 705458
rect 127222 705222 162986 705458
rect 163222 705222 198986 705458
rect 199222 705222 234986 705458
rect 235222 705222 270986 705458
rect 271222 705222 306986 705458
rect 307222 705222 342986 705458
rect 343222 705222 378986 705458
rect 379222 705222 414986 705458
rect 415222 705222 450986 705458
rect 451222 705222 486986 705458
rect 487222 705222 522986 705458
rect 523222 705222 558986 705458
rect 559222 705222 586442 705458
rect 586678 705222 586860 705458
rect -2936 705200 586860 705222
rect -2936 705198 -2336 705200
rect 18804 705198 19404 705200
rect 54804 705198 55404 705200
rect 90804 705198 91404 705200
rect 126804 705198 127404 705200
rect 162804 705198 163404 705200
rect 198804 705198 199404 705200
rect 234804 705198 235404 705200
rect 270804 705198 271404 705200
rect 306804 705198 307404 705200
rect 342804 705198 343404 705200
rect 378804 705198 379404 705200
rect 414804 705198 415404 705200
rect 450804 705198 451404 705200
rect 486804 705198 487404 705200
rect 522804 705198 523404 705200
rect 558804 705198 559404 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2936 686454 586860 686476
rect -2936 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586860 686454
rect -2936 686134 586860 686218
rect -2936 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586860 686134
rect -2936 685876 586860 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -2936 668476 -2336 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586260 668476 586860 668478
rect -2936 668454 586860 668476
rect -2936 668218 -2754 668454
rect -2518 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586442 668454
rect 586678 668218 586860 668454
rect -2936 668134 586860 668218
rect -2936 667898 -2754 668134
rect -2518 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586442 668134
rect 586678 667898 586860 668134
rect -2936 667876 586860 667898
rect -2936 667874 -2336 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586260 667874 586860 667876
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 108804 650476 109404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 216804 650476 217404 650478
rect 252804 650476 253404 650478
rect 288804 650476 289404 650478
rect 324804 650476 325404 650478
rect 360804 650476 361404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 468804 650476 469404 650478
rect 504804 650476 505404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2936 650454 586860 650476
rect -2936 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 324986 650454
rect 325222 650218 360986 650454
rect 361222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586860 650454
rect -2936 650134 586860 650218
rect -2936 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 324986 650134
rect 325222 649898 360986 650134
rect 361222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586860 650134
rect -2936 649876 586860 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 108804 649874 109404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 216804 649874 217404 649876
rect 252804 649874 253404 649876
rect 288804 649874 289404 649876
rect 324804 649874 325404 649876
rect 360804 649874 361404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 468804 649874 469404 649876
rect 504804 649874 505404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -2936 632476 -2336 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 90804 632476 91404 632478
rect 126804 632476 127404 632478
rect 162804 632476 163404 632478
rect 198804 632476 199404 632478
rect 234804 632476 235404 632478
rect 270804 632476 271404 632478
rect 306804 632476 307404 632478
rect 342804 632476 343404 632478
rect 378804 632476 379404 632478
rect 414804 632476 415404 632478
rect 450804 632476 451404 632478
rect 486804 632476 487404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586260 632476 586860 632478
rect -2936 632454 586860 632476
rect -2936 632218 -2754 632454
rect -2518 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 90986 632454
rect 91222 632218 126986 632454
rect 127222 632218 162986 632454
rect 163222 632218 198986 632454
rect 199222 632218 234986 632454
rect 235222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 342986 632454
rect 343222 632218 378986 632454
rect 379222 632218 414986 632454
rect 415222 632218 450986 632454
rect 451222 632218 486986 632454
rect 487222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586442 632454
rect 586678 632218 586860 632454
rect -2936 632134 586860 632218
rect -2936 631898 -2754 632134
rect -2518 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 90986 632134
rect 91222 631898 126986 632134
rect 127222 631898 162986 632134
rect 163222 631898 198986 632134
rect 199222 631898 234986 632134
rect 235222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 342986 632134
rect 343222 631898 378986 632134
rect 379222 631898 414986 632134
rect 415222 631898 450986 632134
rect 451222 631898 486986 632134
rect 487222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586442 632134
rect 586678 631898 586860 632134
rect -2936 631876 586860 631898
rect -2936 631874 -2336 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 90804 631874 91404 631876
rect 126804 631874 127404 631876
rect 162804 631874 163404 631876
rect 198804 631874 199404 631876
rect 234804 631874 235404 631876
rect 270804 631874 271404 631876
rect 306804 631874 307404 631876
rect 342804 631874 343404 631876
rect 378804 631874 379404 631876
rect 414804 631874 415404 631876
rect 450804 631874 451404 631876
rect 486804 631874 487404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586260 631874 586860 631876
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 72804 614476 73404 614478
rect 108804 614476 109404 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 216804 614476 217404 614478
rect 252804 614476 253404 614478
rect 288804 614476 289404 614478
rect 324804 614476 325404 614478
rect 360804 614476 361404 614478
rect 396804 614476 397404 614478
rect 432804 614476 433404 614478
rect 468804 614476 469404 614478
rect 504804 614476 505404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2936 614454 586860 614476
rect -2936 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 72986 614454
rect 73222 614218 108986 614454
rect 109222 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 216986 614454
rect 217222 614218 252986 614454
rect 253222 614218 288986 614454
rect 289222 614218 324986 614454
rect 325222 614218 360986 614454
rect 361222 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 468986 614454
rect 469222 614218 504986 614454
rect 505222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586860 614454
rect -2936 614134 586860 614218
rect -2936 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 72986 614134
rect 73222 613898 108986 614134
rect 109222 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 216986 614134
rect 217222 613898 252986 614134
rect 253222 613898 288986 614134
rect 289222 613898 324986 614134
rect 325222 613898 360986 614134
rect 361222 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 468986 614134
rect 469222 613898 504986 614134
rect 505222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586860 614134
rect -2936 613876 586860 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 72804 613874 73404 613876
rect 108804 613874 109404 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 216804 613874 217404 613876
rect 252804 613874 253404 613876
rect 288804 613874 289404 613876
rect 324804 613874 325404 613876
rect 360804 613874 361404 613876
rect 396804 613874 397404 613876
rect 432804 613874 433404 613876
rect 468804 613874 469404 613876
rect 504804 613874 505404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -2936 596476 -2336 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 90804 596476 91404 596478
rect 126804 596476 127404 596478
rect 162804 596476 163404 596478
rect 198804 596476 199404 596478
rect 234804 596476 235404 596478
rect 270804 596476 271404 596478
rect 306804 596476 307404 596478
rect 342804 596476 343404 596478
rect 378804 596476 379404 596478
rect 414804 596476 415404 596478
rect 450804 596476 451404 596478
rect 486804 596476 487404 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586260 596476 586860 596478
rect -2936 596454 586860 596476
rect -2936 596218 -2754 596454
rect -2518 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 90986 596454
rect 91222 596218 126986 596454
rect 127222 596218 162986 596454
rect 163222 596218 198986 596454
rect 199222 596218 234986 596454
rect 235222 596218 270986 596454
rect 271222 596218 306986 596454
rect 307222 596218 342986 596454
rect 343222 596218 378986 596454
rect 379222 596218 414986 596454
rect 415222 596218 450986 596454
rect 451222 596218 486986 596454
rect 487222 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586442 596454
rect 586678 596218 586860 596454
rect -2936 596134 586860 596218
rect -2936 595898 -2754 596134
rect -2518 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 90986 596134
rect 91222 595898 126986 596134
rect 127222 595898 162986 596134
rect 163222 595898 198986 596134
rect 199222 595898 234986 596134
rect 235222 595898 270986 596134
rect 271222 595898 306986 596134
rect 307222 595898 342986 596134
rect 343222 595898 378986 596134
rect 379222 595898 414986 596134
rect 415222 595898 450986 596134
rect 451222 595898 486986 596134
rect 487222 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586442 596134
rect 586678 595898 586860 596134
rect -2936 595876 586860 595898
rect -2936 595874 -2336 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 90804 595874 91404 595876
rect 126804 595874 127404 595876
rect 162804 595874 163404 595876
rect 198804 595874 199404 595876
rect 234804 595874 235404 595876
rect 270804 595874 271404 595876
rect 306804 595874 307404 595876
rect 342804 595874 343404 595876
rect 378804 595874 379404 595876
rect 414804 595874 415404 595876
rect 450804 595874 451404 595876
rect 486804 595874 487404 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586260 595874 586860 595876
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 47088 578476 47408 578478
rect 77808 578476 78128 578478
rect 108528 578476 108848 578478
rect 139248 578476 139568 578478
rect 169968 578476 170288 578478
rect 200688 578476 201008 578478
rect 231408 578476 231728 578478
rect 262128 578476 262448 578478
rect 288804 578476 289404 578478
rect 339216 578476 339536 578478
rect 369936 578476 370256 578478
rect 400656 578476 400976 578478
rect 431376 578476 431696 578478
rect 462096 578476 462416 578478
rect 492816 578476 493136 578478
rect 523536 578476 523856 578478
rect 554256 578476 554576 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2936 578454 586860 578476
rect -2936 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 47130 578454
rect 47366 578218 77850 578454
rect 78086 578218 108570 578454
rect 108806 578218 139290 578454
rect 139526 578218 170010 578454
rect 170246 578218 200730 578454
rect 200966 578218 231450 578454
rect 231686 578218 262170 578454
rect 262406 578218 288986 578454
rect 289222 578218 339258 578454
rect 339494 578218 369978 578454
rect 370214 578218 400698 578454
rect 400934 578218 431418 578454
rect 431654 578218 462138 578454
rect 462374 578218 492858 578454
rect 493094 578218 523578 578454
rect 523814 578218 554298 578454
rect 554534 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586860 578454
rect -2936 578134 586860 578218
rect -2936 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 47130 578134
rect 47366 577898 77850 578134
rect 78086 577898 108570 578134
rect 108806 577898 139290 578134
rect 139526 577898 170010 578134
rect 170246 577898 200730 578134
rect 200966 577898 231450 578134
rect 231686 577898 262170 578134
rect 262406 577898 288986 578134
rect 289222 577898 339258 578134
rect 339494 577898 369978 578134
rect 370214 577898 400698 578134
rect 400934 577898 431418 578134
rect 431654 577898 462138 578134
rect 462374 577898 492858 578134
rect 493094 577898 523578 578134
rect 523814 577898 554298 578134
rect 554534 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586860 578134
rect -2936 577876 586860 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 47088 577874 47408 577876
rect 77808 577874 78128 577876
rect 108528 577874 108848 577876
rect 139248 577874 139568 577876
rect 169968 577874 170288 577876
rect 200688 577874 201008 577876
rect 231408 577874 231728 577876
rect 262128 577874 262448 577876
rect 288804 577874 289404 577876
rect 339216 577874 339536 577876
rect 369936 577874 370256 577876
rect 400656 577874 400976 577876
rect 431376 577874 431696 577876
rect 462096 577874 462416 577876
rect 492816 577874 493136 577876
rect 523536 577874 523856 577876
rect 554256 577874 554576 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -2936 560476 -2336 560478
rect 18804 560476 19404 560478
rect 31728 560476 32048 560478
rect 62448 560476 62768 560478
rect 93168 560476 93488 560478
rect 123888 560476 124208 560478
rect 154608 560476 154928 560478
rect 185328 560476 185648 560478
rect 216048 560476 216368 560478
rect 246768 560476 247088 560478
rect 270804 560476 271404 560478
rect 306804 560476 307404 560478
rect 323856 560476 324176 560478
rect 354576 560476 354896 560478
rect 385296 560476 385616 560478
rect 416016 560476 416336 560478
rect 446736 560476 447056 560478
rect 477456 560476 477776 560478
rect 508176 560476 508496 560478
rect 538896 560476 539216 560478
rect 586260 560476 586860 560478
rect -2936 560454 586860 560476
rect -2936 560218 -2754 560454
rect -2518 560218 18986 560454
rect 19222 560218 31770 560454
rect 32006 560218 62490 560454
rect 62726 560218 93210 560454
rect 93446 560218 123930 560454
rect 124166 560218 154650 560454
rect 154886 560218 185370 560454
rect 185606 560218 216090 560454
rect 216326 560218 246810 560454
rect 247046 560218 270986 560454
rect 271222 560218 306986 560454
rect 307222 560218 323898 560454
rect 324134 560218 354618 560454
rect 354854 560218 385338 560454
rect 385574 560218 416058 560454
rect 416294 560218 446778 560454
rect 447014 560218 477498 560454
rect 477734 560218 508218 560454
rect 508454 560218 538938 560454
rect 539174 560218 586442 560454
rect 586678 560218 586860 560454
rect -2936 560134 586860 560218
rect -2936 559898 -2754 560134
rect -2518 559898 18986 560134
rect 19222 559898 31770 560134
rect 32006 559898 62490 560134
rect 62726 559898 93210 560134
rect 93446 559898 123930 560134
rect 124166 559898 154650 560134
rect 154886 559898 185370 560134
rect 185606 559898 216090 560134
rect 216326 559898 246810 560134
rect 247046 559898 270986 560134
rect 271222 559898 306986 560134
rect 307222 559898 323898 560134
rect 324134 559898 354618 560134
rect 354854 559898 385338 560134
rect 385574 559898 416058 560134
rect 416294 559898 446778 560134
rect 447014 559898 477498 560134
rect 477734 559898 508218 560134
rect 508454 559898 538938 560134
rect 539174 559898 586442 560134
rect 586678 559898 586860 560134
rect -2936 559876 586860 559898
rect -2936 559874 -2336 559876
rect 18804 559874 19404 559876
rect 31728 559874 32048 559876
rect 62448 559874 62768 559876
rect 93168 559874 93488 559876
rect 123888 559874 124208 559876
rect 154608 559874 154928 559876
rect 185328 559874 185648 559876
rect 216048 559874 216368 559876
rect 246768 559874 247088 559876
rect 270804 559874 271404 559876
rect 306804 559874 307404 559876
rect 323856 559874 324176 559876
rect 354576 559874 354896 559876
rect 385296 559874 385616 559876
rect 416016 559874 416336 559876
rect 446736 559874 447056 559876
rect 477456 559874 477776 559876
rect 508176 559874 508496 559876
rect 538896 559874 539216 559876
rect 586260 559874 586860 559876
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 47088 542476 47408 542478
rect 77808 542476 78128 542478
rect 108528 542476 108848 542478
rect 139248 542476 139568 542478
rect 169968 542476 170288 542478
rect 200688 542476 201008 542478
rect 231408 542476 231728 542478
rect 262128 542476 262448 542478
rect 288804 542476 289404 542478
rect 339216 542476 339536 542478
rect 369936 542476 370256 542478
rect 400656 542476 400976 542478
rect 431376 542476 431696 542478
rect 462096 542476 462416 542478
rect 492816 542476 493136 542478
rect 523536 542476 523856 542478
rect 554256 542476 554576 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2936 542454 586860 542476
rect -2936 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 47130 542454
rect 47366 542218 77850 542454
rect 78086 542218 108570 542454
rect 108806 542218 139290 542454
rect 139526 542218 170010 542454
rect 170246 542218 200730 542454
rect 200966 542218 231450 542454
rect 231686 542218 262170 542454
rect 262406 542218 288986 542454
rect 289222 542218 339258 542454
rect 339494 542218 369978 542454
rect 370214 542218 400698 542454
rect 400934 542218 431418 542454
rect 431654 542218 462138 542454
rect 462374 542218 492858 542454
rect 493094 542218 523578 542454
rect 523814 542218 554298 542454
rect 554534 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586860 542454
rect -2936 542134 586860 542218
rect -2936 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 47130 542134
rect 47366 541898 77850 542134
rect 78086 541898 108570 542134
rect 108806 541898 139290 542134
rect 139526 541898 170010 542134
rect 170246 541898 200730 542134
rect 200966 541898 231450 542134
rect 231686 541898 262170 542134
rect 262406 541898 288986 542134
rect 289222 541898 339258 542134
rect 339494 541898 369978 542134
rect 370214 541898 400698 542134
rect 400934 541898 431418 542134
rect 431654 541898 462138 542134
rect 462374 541898 492858 542134
rect 493094 541898 523578 542134
rect 523814 541898 554298 542134
rect 554534 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586860 542134
rect -2936 541876 586860 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 47088 541874 47408 541876
rect 77808 541874 78128 541876
rect 108528 541874 108848 541876
rect 139248 541874 139568 541876
rect 169968 541874 170288 541876
rect 200688 541874 201008 541876
rect 231408 541874 231728 541876
rect 262128 541874 262448 541876
rect 288804 541874 289404 541876
rect 339216 541874 339536 541876
rect 369936 541874 370256 541876
rect 400656 541874 400976 541876
rect 431376 541874 431696 541876
rect 462096 541874 462416 541876
rect 492816 541874 493136 541876
rect 523536 541874 523856 541876
rect 554256 541874 554576 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -2936 524476 -2336 524478
rect 18804 524476 19404 524478
rect 31728 524476 32048 524478
rect 62448 524476 62768 524478
rect 93168 524476 93488 524478
rect 123888 524476 124208 524478
rect 154608 524476 154928 524478
rect 185328 524476 185648 524478
rect 216048 524476 216368 524478
rect 246768 524476 247088 524478
rect 270804 524476 271404 524478
rect 306804 524476 307404 524478
rect 323856 524476 324176 524478
rect 354576 524476 354896 524478
rect 385296 524476 385616 524478
rect 416016 524476 416336 524478
rect 446736 524476 447056 524478
rect 477456 524476 477776 524478
rect 508176 524476 508496 524478
rect 538896 524476 539216 524478
rect 586260 524476 586860 524478
rect -2936 524454 586860 524476
rect -2936 524218 -2754 524454
rect -2518 524218 18986 524454
rect 19222 524218 31770 524454
rect 32006 524218 62490 524454
rect 62726 524218 93210 524454
rect 93446 524218 123930 524454
rect 124166 524218 154650 524454
rect 154886 524218 185370 524454
rect 185606 524218 216090 524454
rect 216326 524218 246810 524454
rect 247046 524218 270986 524454
rect 271222 524218 306986 524454
rect 307222 524218 323898 524454
rect 324134 524218 354618 524454
rect 354854 524218 385338 524454
rect 385574 524218 416058 524454
rect 416294 524218 446778 524454
rect 447014 524218 477498 524454
rect 477734 524218 508218 524454
rect 508454 524218 538938 524454
rect 539174 524218 586442 524454
rect 586678 524218 586860 524454
rect -2936 524134 586860 524218
rect -2936 523898 -2754 524134
rect -2518 523898 18986 524134
rect 19222 523898 31770 524134
rect 32006 523898 62490 524134
rect 62726 523898 93210 524134
rect 93446 523898 123930 524134
rect 124166 523898 154650 524134
rect 154886 523898 185370 524134
rect 185606 523898 216090 524134
rect 216326 523898 246810 524134
rect 247046 523898 270986 524134
rect 271222 523898 306986 524134
rect 307222 523898 323898 524134
rect 324134 523898 354618 524134
rect 354854 523898 385338 524134
rect 385574 523898 416058 524134
rect 416294 523898 446778 524134
rect 447014 523898 477498 524134
rect 477734 523898 508218 524134
rect 508454 523898 538938 524134
rect 539174 523898 586442 524134
rect 586678 523898 586860 524134
rect -2936 523876 586860 523898
rect -2936 523874 -2336 523876
rect 18804 523874 19404 523876
rect 31728 523874 32048 523876
rect 62448 523874 62768 523876
rect 93168 523874 93488 523876
rect 123888 523874 124208 523876
rect 154608 523874 154928 523876
rect 185328 523874 185648 523876
rect 216048 523874 216368 523876
rect 246768 523874 247088 523876
rect 270804 523874 271404 523876
rect 306804 523874 307404 523876
rect 323856 523874 324176 523876
rect 354576 523874 354896 523876
rect 385296 523874 385616 523876
rect 416016 523874 416336 523876
rect 446736 523874 447056 523876
rect 477456 523874 477776 523876
rect 508176 523874 508496 523876
rect 538896 523874 539216 523876
rect 586260 523874 586860 523876
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 47088 506476 47408 506478
rect 77808 506476 78128 506478
rect 108528 506476 108848 506478
rect 139248 506476 139568 506478
rect 169968 506476 170288 506478
rect 200688 506476 201008 506478
rect 231408 506476 231728 506478
rect 262128 506476 262448 506478
rect 288804 506476 289404 506478
rect 339216 506476 339536 506478
rect 369936 506476 370256 506478
rect 400656 506476 400976 506478
rect 431376 506476 431696 506478
rect 462096 506476 462416 506478
rect 492816 506476 493136 506478
rect 523536 506476 523856 506478
rect 554256 506476 554576 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2936 506454 586860 506476
rect -2936 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 47130 506454
rect 47366 506218 77850 506454
rect 78086 506218 108570 506454
rect 108806 506218 139290 506454
rect 139526 506218 170010 506454
rect 170246 506218 200730 506454
rect 200966 506218 231450 506454
rect 231686 506218 262170 506454
rect 262406 506218 288986 506454
rect 289222 506218 339258 506454
rect 339494 506218 369978 506454
rect 370214 506218 400698 506454
rect 400934 506218 431418 506454
rect 431654 506218 462138 506454
rect 462374 506218 492858 506454
rect 493094 506218 523578 506454
rect 523814 506218 554298 506454
rect 554534 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586860 506454
rect -2936 506134 586860 506218
rect -2936 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 47130 506134
rect 47366 505898 77850 506134
rect 78086 505898 108570 506134
rect 108806 505898 139290 506134
rect 139526 505898 170010 506134
rect 170246 505898 200730 506134
rect 200966 505898 231450 506134
rect 231686 505898 262170 506134
rect 262406 505898 288986 506134
rect 289222 505898 339258 506134
rect 339494 505898 369978 506134
rect 370214 505898 400698 506134
rect 400934 505898 431418 506134
rect 431654 505898 462138 506134
rect 462374 505898 492858 506134
rect 493094 505898 523578 506134
rect 523814 505898 554298 506134
rect 554534 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586860 506134
rect -2936 505876 586860 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 47088 505874 47408 505876
rect 77808 505874 78128 505876
rect 108528 505874 108848 505876
rect 139248 505874 139568 505876
rect 169968 505874 170288 505876
rect 200688 505874 201008 505876
rect 231408 505874 231728 505876
rect 262128 505874 262448 505876
rect 288804 505874 289404 505876
rect 339216 505874 339536 505876
rect 369936 505874 370256 505876
rect 400656 505874 400976 505876
rect 431376 505874 431696 505876
rect 462096 505874 462416 505876
rect 492816 505874 493136 505876
rect 523536 505874 523856 505876
rect 554256 505874 554576 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -2936 488476 -2336 488478
rect 18804 488476 19404 488478
rect 31728 488476 32048 488478
rect 62448 488476 62768 488478
rect 93168 488476 93488 488478
rect 123888 488476 124208 488478
rect 154608 488476 154928 488478
rect 185328 488476 185648 488478
rect 216048 488476 216368 488478
rect 246768 488476 247088 488478
rect 270804 488476 271404 488478
rect 306804 488476 307404 488478
rect 323856 488476 324176 488478
rect 354576 488476 354896 488478
rect 385296 488476 385616 488478
rect 416016 488476 416336 488478
rect 446736 488476 447056 488478
rect 477456 488476 477776 488478
rect 508176 488476 508496 488478
rect 538896 488476 539216 488478
rect 586260 488476 586860 488478
rect -2936 488454 586860 488476
rect -2936 488218 -2754 488454
rect -2518 488218 18986 488454
rect 19222 488218 31770 488454
rect 32006 488218 62490 488454
rect 62726 488218 93210 488454
rect 93446 488218 123930 488454
rect 124166 488218 154650 488454
rect 154886 488218 185370 488454
rect 185606 488218 216090 488454
rect 216326 488218 246810 488454
rect 247046 488218 270986 488454
rect 271222 488218 306986 488454
rect 307222 488218 323898 488454
rect 324134 488218 354618 488454
rect 354854 488218 385338 488454
rect 385574 488218 416058 488454
rect 416294 488218 446778 488454
rect 447014 488218 477498 488454
rect 477734 488218 508218 488454
rect 508454 488218 538938 488454
rect 539174 488218 586442 488454
rect 586678 488218 586860 488454
rect -2936 488134 586860 488218
rect -2936 487898 -2754 488134
rect -2518 487898 18986 488134
rect 19222 487898 31770 488134
rect 32006 487898 62490 488134
rect 62726 487898 93210 488134
rect 93446 487898 123930 488134
rect 124166 487898 154650 488134
rect 154886 487898 185370 488134
rect 185606 487898 216090 488134
rect 216326 487898 246810 488134
rect 247046 487898 270986 488134
rect 271222 487898 306986 488134
rect 307222 487898 323898 488134
rect 324134 487898 354618 488134
rect 354854 487898 385338 488134
rect 385574 487898 416058 488134
rect 416294 487898 446778 488134
rect 447014 487898 477498 488134
rect 477734 487898 508218 488134
rect 508454 487898 538938 488134
rect 539174 487898 586442 488134
rect 586678 487898 586860 488134
rect -2936 487876 586860 487898
rect -2936 487874 -2336 487876
rect 18804 487874 19404 487876
rect 31728 487874 32048 487876
rect 62448 487874 62768 487876
rect 93168 487874 93488 487876
rect 123888 487874 124208 487876
rect 154608 487874 154928 487876
rect 185328 487874 185648 487876
rect 216048 487874 216368 487876
rect 246768 487874 247088 487876
rect 270804 487874 271404 487876
rect 306804 487874 307404 487876
rect 323856 487874 324176 487876
rect 354576 487874 354896 487876
rect 385296 487874 385616 487876
rect 416016 487874 416336 487876
rect 446736 487874 447056 487876
rect 477456 487874 477776 487876
rect 508176 487874 508496 487876
rect 538896 487874 539216 487876
rect 586260 487874 586860 487876
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 47088 470476 47408 470478
rect 77808 470476 78128 470478
rect 108528 470476 108848 470478
rect 139248 470476 139568 470478
rect 169968 470476 170288 470478
rect 200688 470476 201008 470478
rect 231408 470476 231728 470478
rect 262128 470476 262448 470478
rect 288804 470476 289404 470478
rect 339216 470476 339536 470478
rect 369936 470476 370256 470478
rect 400656 470476 400976 470478
rect 431376 470476 431696 470478
rect 462096 470476 462416 470478
rect 492816 470476 493136 470478
rect 523536 470476 523856 470478
rect 554256 470476 554576 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2936 470454 586860 470476
rect -2936 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 47130 470454
rect 47366 470218 77850 470454
rect 78086 470218 108570 470454
rect 108806 470218 139290 470454
rect 139526 470218 170010 470454
rect 170246 470218 200730 470454
rect 200966 470218 231450 470454
rect 231686 470218 262170 470454
rect 262406 470218 288986 470454
rect 289222 470218 339258 470454
rect 339494 470218 369978 470454
rect 370214 470218 400698 470454
rect 400934 470218 431418 470454
rect 431654 470218 462138 470454
rect 462374 470218 492858 470454
rect 493094 470218 523578 470454
rect 523814 470218 554298 470454
rect 554534 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586860 470454
rect -2936 470134 586860 470218
rect -2936 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 47130 470134
rect 47366 469898 77850 470134
rect 78086 469898 108570 470134
rect 108806 469898 139290 470134
rect 139526 469898 170010 470134
rect 170246 469898 200730 470134
rect 200966 469898 231450 470134
rect 231686 469898 262170 470134
rect 262406 469898 288986 470134
rect 289222 469898 339258 470134
rect 339494 469898 369978 470134
rect 370214 469898 400698 470134
rect 400934 469898 431418 470134
rect 431654 469898 462138 470134
rect 462374 469898 492858 470134
rect 493094 469898 523578 470134
rect 523814 469898 554298 470134
rect 554534 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586860 470134
rect -2936 469876 586860 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 47088 469874 47408 469876
rect 77808 469874 78128 469876
rect 108528 469874 108848 469876
rect 139248 469874 139568 469876
rect 169968 469874 170288 469876
rect 200688 469874 201008 469876
rect 231408 469874 231728 469876
rect 262128 469874 262448 469876
rect 288804 469874 289404 469876
rect 339216 469874 339536 469876
rect 369936 469874 370256 469876
rect 400656 469874 400976 469876
rect 431376 469874 431696 469876
rect 462096 469874 462416 469876
rect 492816 469874 493136 469876
rect 523536 469874 523856 469876
rect 554256 469874 554576 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -2936 452476 -2336 452478
rect 18804 452476 19404 452478
rect 31728 452476 32048 452478
rect 62448 452476 62768 452478
rect 93168 452476 93488 452478
rect 123888 452476 124208 452478
rect 154608 452476 154928 452478
rect 185328 452476 185648 452478
rect 216048 452476 216368 452478
rect 246768 452476 247088 452478
rect 270804 452476 271404 452478
rect 306804 452476 307404 452478
rect 323856 452476 324176 452478
rect 354576 452476 354896 452478
rect 385296 452476 385616 452478
rect 416016 452476 416336 452478
rect 446736 452476 447056 452478
rect 477456 452476 477776 452478
rect 508176 452476 508496 452478
rect 538896 452476 539216 452478
rect 586260 452476 586860 452478
rect -2936 452454 586860 452476
rect -2936 452218 -2754 452454
rect -2518 452218 18986 452454
rect 19222 452218 31770 452454
rect 32006 452218 62490 452454
rect 62726 452218 93210 452454
rect 93446 452218 123930 452454
rect 124166 452218 154650 452454
rect 154886 452218 185370 452454
rect 185606 452218 216090 452454
rect 216326 452218 246810 452454
rect 247046 452218 270986 452454
rect 271222 452218 306986 452454
rect 307222 452218 323898 452454
rect 324134 452218 354618 452454
rect 354854 452218 385338 452454
rect 385574 452218 416058 452454
rect 416294 452218 446778 452454
rect 447014 452218 477498 452454
rect 477734 452218 508218 452454
rect 508454 452218 538938 452454
rect 539174 452218 586442 452454
rect 586678 452218 586860 452454
rect -2936 452134 586860 452218
rect -2936 451898 -2754 452134
rect -2518 451898 18986 452134
rect 19222 451898 31770 452134
rect 32006 451898 62490 452134
rect 62726 451898 93210 452134
rect 93446 451898 123930 452134
rect 124166 451898 154650 452134
rect 154886 451898 185370 452134
rect 185606 451898 216090 452134
rect 216326 451898 246810 452134
rect 247046 451898 270986 452134
rect 271222 451898 306986 452134
rect 307222 451898 323898 452134
rect 324134 451898 354618 452134
rect 354854 451898 385338 452134
rect 385574 451898 416058 452134
rect 416294 451898 446778 452134
rect 447014 451898 477498 452134
rect 477734 451898 508218 452134
rect 508454 451898 538938 452134
rect 539174 451898 586442 452134
rect 586678 451898 586860 452134
rect -2936 451876 586860 451898
rect -2936 451874 -2336 451876
rect 18804 451874 19404 451876
rect 31728 451874 32048 451876
rect 62448 451874 62768 451876
rect 93168 451874 93488 451876
rect 123888 451874 124208 451876
rect 154608 451874 154928 451876
rect 185328 451874 185648 451876
rect 216048 451874 216368 451876
rect 246768 451874 247088 451876
rect 270804 451874 271404 451876
rect 306804 451874 307404 451876
rect 323856 451874 324176 451876
rect 354576 451874 354896 451876
rect 385296 451874 385616 451876
rect 416016 451874 416336 451876
rect 446736 451874 447056 451876
rect 477456 451874 477776 451876
rect 508176 451874 508496 451876
rect 538896 451874 539216 451876
rect 586260 451874 586860 451876
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 47088 434476 47408 434478
rect 77808 434476 78128 434478
rect 108528 434476 108848 434478
rect 139248 434476 139568 434478
rect 169968 434476 170288 434478
rect 200688 434476 201008 434478
rect 231408 434476 231728 434478
rect 262128 434476 262448 434478
rect 288804 434476 289404 434478
rect 339216 434476 339536 434478
rect 369936 434476 370256 434478
rect 400656 434476 400976 434478
rect 431376 434476 431696 434478
rect 462096 434476 462416 434478
rect 492816 434476 493136 434478
rect 523536 434476 523856 434478
rect 554256 434476 554576 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2936 434454 586860 434476
rect -2936 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 47130 434454
rect 47366 434218 77850 434454
rect 78086 434218 108570 434454
rect 108806 434218 139290 434454
rect 139526 434218 170010 434454
rect 170246 434218 200730 434454
rect 200966 434218 231450 434454
rect 231686 434218 262170 434454
rect 262406 434218 288986 434454
rect 289222 434218 339258 434454
rect 339494 434218 369978 434454
rect 370214 434218 400698 434454
rect 400934 434218 431418 434454
rect 431654 434218 462138 434454
rect 462374 434218 492858 434454
rect 493094 434218 523578 434454
rect 523814 434218 554298 434454
rect 554534 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586860 434454
rect -2936 434134 586860 434218
rect -2936 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 47130 434134
rect 47366 433898 77850 434134
rect 78086 433898 108570 434134
rect 108806 433898 139290 434134
rect 139526 433898 170010 434134
rect 170246 433898 200730 434134
rect 200966 433898 231450 434134
rect 231686 433898 262170 434134
rect 262406 433898 288986 434134
rect 289222 433898 339258 434134
rect 339494 433898 369978 434134
rect 370214 433898 400698 434134
rect 400934 433898 431418 434134
rect 431654 433898 462138 434134
rect 462374 433898 492858 434134
rect 493094 433898 523578 434134
rect 523814 433898 554298 434134
rect 554534 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586860 434134
rect -2936 433876 586860 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 47088 433874 47408 433876
rect 77808 433874 78128 433876
rect 108528 433874 108848 433876
rect 139248 433874 139568 433876
rect 169968 433874 170288 433876
rect 200688 433874 201008 433876
rect 231408 433874 231728 433876
rect 262128 433874 262448 433876
rect 288804 433874 289404 433876
rect 339216 433874 339536 433876
rect 369936 433874 370256 433876
rect 400656 433874 400976 433876
rect 431376 433874 431696 433876
rect 462096 433874 462416 433876
rect 492816 433874 493136 433876
rect 523536 433874 523856 433876
rect 554256 433874 554576 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -2936 416476 -2336 416478
rect 18804 416476 19404 416478
rect 31728 416476 32048 416478
rect 62448 416476 62768 416478
rect 93168 416476 93488 416478
rect 123888 416476 124208 416478
rect 154608 416476 154928 416478
rect 185328 416476 185648 416478
rect 216048 416476 216368 416478
rect 246768 416476 247088 416478
rect 270804 416476 271404 416478
rect 306804 416476 307404 416478
rect 323856 416476 324176 416478
rect 354576 416476 354896 416478
rect 385296 416476 385616 416478
rect 416016 416476 416336 416478
rect 446736 416476 447056 416478
rect 477456 416476 477776 416478
rect 508176 416476 508496 416478
rect 538896 416476 539216 416478
rect 586260 416476 586860 416478
rect -2936 416454 586860 416476
rect -2936 416218 -2754 416454
rect -2518 416218 18986 416454
rect 19222 416218 31770 416454
rect 32006 416218 62490 416454
rect 62726 416218 93210 416454
rect 93446 416218 123930 416454
rect 124166 416218 154650 416454
rect 154886 416218 185370 416454
rect 185606 416218 216090 416454
rect 216326 416218 246810 416454
rect 247046 416218 270986 416454
rect 271222 416218 306986 416454
rect 307222 416218 323898 416454
rect 324134 416218 354618 416454
rect 354854 416218 385338 416454
rect 385574 416218 416058 416454
rect 416294 416218 446778 416454
rect 447014 416218 477498 416454
rect 477734 416218 508218 416454
rect 508454 416218 538938 416454
rect 539174 416218 586442 416454
rect 586678 416218 586860 416454
rect -2936 416134 586860 416218
rect -2936 415898 -2754 416134
rect -2518 415898 18986 416134
rect 19222 415898 31770 416134
rect 32006 415898 62490 416134
rect 62726 415898 93210 416134
rect 93446 415898 123930 416134
rect 124166 415898 154650 416134
rect 154886 415898 185370 416134
rect 185606 415898 216090 416134
rect 216326 415898 246810 416134
rect 247046 415898 270986 416134
rect 271222 415898 306986 416134
rect 307222 415898 323898 416134
rect 324134 415898 354618 416134
rect 354854 415898 385338 416134
rect 385574 415898 416058 416134
rect 416294 415898 446778 416134
rect 447014 415898 477498 416134
rect 477734 415898 508218 416134
rect 508454 415898 538938 416134
rect 539174 415898 586442 416134
rect 586678 415898 586860 416134
rect -2936 415876 586860 415898
rect -2936 415874 -2336 415876
rect 18804 415874 19404 415876
rect 31728 415874 32048 415876
rect 62448 415874 62768 415876
rect 93168 415874 93488 415876
rect 123888 415874 124208 415876
rect 154608 415874 154928 415876
rect 185328 415874 185648 415876
rect 216048 415874 216368 415876
rect 246768 415874 247088 415876
rect 270804 415874 271404 415876
rect 306804 415874 307404 415876
rect 323856 415874 324176 415876
rect 354576 415874 354896 415876
rect 385296 415874 385616 415876
rect 416016 415874 416336 415876
rect 446736 415874 447056 415876
rect 477456 415874 477776 415876
rect 508176 415874 508496 415876
rect 538896 415874 539216 415876
rect 586260 415874 586860 415876
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 47088 398476 47408 398478
rect 77808 398476 78128 398478
rect 108528 398476 108848 398478
rect 139248 398476 139568 398478
rect 169968 398476 170288 398478
rect 200688 398476 201008 398478
rect 231408 398476 231728 398478
rect 262128 398476 262448 398478
rect 288804 398476 289404 398478
rect 339216 398476 339536 398478
rect 369936 398476 370256 398478
rect 400656 398476 400976 398478
rect 431376 398476 431696 398478
rect 462096 398476 462416 398478
rect 492816 398476 493136 398478
rect 523536 398476 523856 398478
rect 554256 398476 554576 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2936 398454 586860 398476
rect -2936 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 47130 398454
rect 47366 398218 77850 398454
rect 78086 398218 108570 398454
rect 108806 398218 139290 398454
rect 139526 398218 170010 398454
rect 170246 398218 200730 398454
rect 200966 398218 231450 398454
rect 231686 398218 262170 398454
rect 262406 398218 288986 398454
rect 289222 398218 339258 398454
rect 339494 398218 369978 398454
rect 370214 398218 400698 398454
rect 400934 398218 431418 398454
rect 431654 398218 462138 398454
rect 462374 398218 492858 398454
rect 493094 398218 523578 398454
rect 523814 398218 554298 398454
rect 554534 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586860 398454
rect -2936 398134 586860 398218
rect -2936 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 47130 398134
rect 47366 397898 77850 398134
rect 78086 397898 108570 398134
rect 108806 397898 139290 398134
rect 139526 397898 170010 398134
rect 170246 397898 200730 398134
rect 200966 397898 231450 398134
rect 231686 397898 262170 398134
rect 262406 397898 288986 398134
rect 289222 397898 339258 398134
rect 339494 397898 369978 398134
rect 370214 397898 400698 398134
rect 400934 397898 431418 398134
rect 431654 397898 462138 398134
rect 462374 397898 492858 398134
rect 493094 397898 523578 398134
rect 523814 397898 554298 398134
rect 554534 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586860 398134
rect -2936 397876 586860 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 47088 397874 47408 397876
rect 77808 397874 78128 397876
rect 108528 397874 108848 397876
rect 139248 397874 139568 397876
rect 169968 397874 170288 397876
rect 200688 397874 201008 397876
rect 231408 397874 231728 397876
rect 262128 397874 262448 397876
rect 288804 397874 289404 397876
rect 339216 397874 339536 397876
rect 369936 397874 370256 397876
rect 400656 397874 400976 397876
rect 431376 397874 431696 397876
rect 462096 397874 462416 397876
rect 492816 397874 493136 397876
rect 523536 397874 523856 397876
rect 554256 397874 554576 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -2936 380476 -2336 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 90804 380476 91404 380478
rect 126804 380476 127404 380478
rect 162804 380476 163404 380478
rect 198804 380476 199404 380478
rect 234804 380476 235404 380478
rect 270804 380476 271404 380478
rect 306804 380476 307404 380478
rect 342804 380476 343404 380478
rect 378804 380476 379404 380478
rect 414804 380476 415404 380478
rect 450804 380476 451404 380478
rect 486804 380476 487404 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586260 380476 586860 380478
rect -2936 380454 586860 380476
rect -2936 380218 -2754 380454
rect -2518 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 90986 380454
rect 91222 380218 126986 380454
rect 127222 380218 162986 380454
rect 163222 380218 198986 380454
rect 199222 380218 234986 380454
rect 235222 380218 270986 380454
rect 271222 380218 306986 380454
rect 307222 380218 342986 380454
rect 343222 380218 378986 380454
rect 379222 380218 414986 380454
rect 415222 380218 450986 380454
rect 451222 380218 486986 380454
rect 487222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586442 380454
rect 586678 380218 586860 380454
rect -2936 380134 586860 380218
rect -2936 379898 -2754 380134
rect -2518 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 90986 380134
rect 91222 379898 126986 380134
rect 127222 379898 162986 380134
rect 163222 379898 198986 380134
rect 199222 379898 234986 380134
rect 235222 379898 270986 380134
rect 271222 379898 306986 380134
rect 307222 379898 342986 380134
rect 343222 379898 378986 380134
rect 379222 379898 414986 380134
rect 415222 379898 450986 380134
rect 451222 379898 486986 380134
rect 487222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586442 380134
rect 586678 379898 586860 380134
rect -2936 379876 586860 379898
rect -2936 379874 -2336 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 90804 379874 91404 379876
rect 126804 379874 127404 379876
rect 162804 379874 163404 379876
rect 198804 379874 199404 379876
rect 234804 379874 235404 379876
rect 270804 379874 271404 379876
rect 306804 379874 307404 379876
rect 342804 379874 343404 379876
rect 378804 379874 379404 379876
rect 414804 379874 415404 379876
rect 450804 379874 451404 379876
rect 486804 379874 487404 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586260 379874 586860 379876
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 72804 362476 73404 362478
rect 108804 362476 109404 362478
rect 144804 362476 145404 362478
rect 180804 362476 181404 362478
rect 216804 362476 217404 362478
rect 252804 362476 253404 362478
rect 288804 362476 289404 362478
rect 324804 362476 325404 362478
rect 360804 362476 361404 362478
rect 396804 362476 397404 362478
rect 432804 362476 433404 362478
rect 468804 362476 469404 362478
rect 504804 362476 505404 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2936 362454 586860 362476
rect -2936 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 72986 362454
rect 73222 362218 108986 362454
rect 109222 362218 144986 362454
rect 145222 362218 180986 362454
rect 181222 362218 216986 362454
rect 217222 362218 252986 362454
rect 253222 362218 288986 362454
rect 289222 362218 324986 362454
rect 325222 362218 360986 362454
rect 361222 362218 396986 362454
rect 397222 362218 432986 362454
rect 433222 362218 468986 362454
rect 469222 362218 504986 362454
rect 505222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586860 362454
rect -2936 362134 586860 362218
rect -2936 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 72986 362134
rect 73222 361898 108986 362134
rect 109222 361898 144986 362134
rect 145222 361898 180986 362134
rect 181222 361898 216986 362134
rect 217222 361898 252986 362134
rect 253222 361898 288986 362134
rect 289222 361898 324986 362134
rect 325222 361898 360986 362134
rect 361222 361898 396986 362134
rect 397222 361898 432986 362134
rect 433222 361898 468986 362134
rect 469222 361898 504986 362134
rect 505222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586860 362134
rect -2936 361876 586860 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 72804 361874 73404 361876
rect 108804 361874 109404 361876
rect 144804 361874 145404 361876
rect 180804 361874 181404 361876
rect 216804 361874 217404 361876
rect 252804 361874 253404 361876
rect 288804 361874 289404 361876
rect 324804 361874 325404 361876
rect 360804 361874 361404 361876
rect 396804 361874 397404 361876
rect 432804 361874 433404 361876
rect 468804 361874 469404 361876
rect 504804 361874 505404 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -2936 344476 -2336 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 90804 344476 91404 344478
rect 126804 344476 127404 344478
rect 162804 344476 163404 344478
rect 198804 344476 199404 344478
rect 234804 344476 235404 344478
rect 292112 344476 292432 344478
rect 342804 344476 343404 344478
rect 378804 344476 379404 344478
rect 414804 344476 415404 344478
rect 450804 344476 451404 344478
rect 486804 344476 487404 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586260 344476 586860 344478
rect -2936 344454 586860 344476
rect -2936 344218 -2754 344454
rect -2518 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 90986 344454
rect 91222 344218 126986 344454
rect 127222 344218 162986 344454
rect 163222 344218 198986 344454
rect 199222 344218 234986 344454
rect 235222 344218 292154 344454
rect 292390 344218 342986 344454
rect 343222 344218 378986 344454
rect 379222 344218 414986 344454
rect 415222 344218 450986 344454
rect 451222 344218 486986 344454
rect 487222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586442 344454
rect 586678 344218 586860 344454
rect -2936 344134 586860 344218
rect -2936 343898 -2754 344134
rect -2518 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 90986 344134
rect 91222 343898 126986 344134
rect 127222 343898 162986 344134
rect 163222 343898 198986 344134
rect 199222 343898 234986 344134
rect 235222 343898 292154 344134
rect 292390 343898 342986 344134
rect 343222 343898 378986 344134
rect 379222 343898 414986 344134
rect 415222 343898 450986 344134
rect 451222 343898 486986 344134
rect 487222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586442 344134
rect 586678 343898 586860 344134
rect -2936 343876 586860 343898
rect -2936 343874 -2336 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 90804 343874 91404 343876
rect 126804 343874 127404 343876
rect 162804 343874 163404 343876
rect 198804 343874 199404 343876
rect 234804 343874 235404 343876
rect 292112 343874 292432 343876
rect 342804 343874 343404 343876
rect 378804 343874 379404 343876
rect 414804 343874 415404 343876
rect 450804 343874 451404 343876
rect 486804 343874 487404 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586260 343874 586860 343876
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 72804 326476 73404 326478
rect 108804 326476 109404 326478
rect 144804 326476 145404 326478
rect 180804 326476 181404 326478
rect 216804 326476 217404 326478
rect 252804 326476 253404 326478
rect 276752 326476 277072 326478
rect 307472 326476 307792 326478
rect 324804 326476 325404 326478
rect 360804 326476 361404 326478
rect 396804 326476 397404 326478
rect 432804 326476 433404 326478
rect 468804 326476 469404 326478
rect 504804 326476 505404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2936 326454 586860 326476
rect -2936 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 72986 326454
rect 73222 326218 108986 326454
rect 109222 326218 144986 326454
rect 145222 326218 180986 326454
rect 181222 326218 216986 326454
rect 217222 326218 252986 326454
rect 253222 326218 276794 326454
rect 277030 326218 307514 326454
rect 307750 326218 324986 326454
rect 325222 326218 360986 326454
rect 361222 326218 396986 326454
rect 397222 326218 432986 326454
rect 433222 326218 468986 326454
rect 469222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586860 326454
rect -2936 326134 586860 326218
rect -2936 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 72986 326134
rect 73222 325898 108986 326134
rect 109222 325898 144986 326134
rect 145222 325898 180986 326134
rect 181222 325898 216986 326134
rect 217222 325898 252986 326134
rect 253222 325898 276794 326134
rect 277030 325898 307514 326134
rect 307750 325898 324986 326134
rect 325222 325898 360986 326134
rect 361222 325898 396986 326134
rect 397222 325898 432986 326134
rect 433222 325898 468986 326134
rect 469222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586860 326134
rect -2936 325876 586860 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 72804 325874 73404 325876
rect 108804 325874 109404 325876
rect 144804 325874 145404 325876
rect 180804 325874 181404 325876
rect 216804 325874 217404 325876
rect 252804 325874 253404 325876
rect 276752 325874 277072 325876
rect 307472 325874 307792 325876
rect 324804 325874 325404 325876
rect 360804 325874 361404 325876
rect 396804 325874 397404 325876
rect 432804 325874 433404 325876
rect 468804 325874 469404 325876
rect 504804 325874 505404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -2936 308476 -2336 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 90804 308476 91404 308478
rect 126804 308476 127404 308478
rect 162804 308476 163404 308478
rect 198804 308476 199404 308478
rect 234804 308476 235404 308478
rect 270804 308476 271404 308478
rect 306804 308476 307404 308478
rect 342804 308476 343404 308478
rect 378804 308476 379404 308478
rect 414804 308476 415404 308478
rect 450804 308476 451404 308478
rect 486804 308476 487404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586260 308476 586860 308478
rect -2936 308454 586860 308476
rect -2936 308218 -2754 308454
rect -2518 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 90986 308454
rect 91222 308218 126986 308454
rect 127222 308218 162986 308454
rect 163222 308218 198986 308454
rect 199222 308218 234986 308454
rect 235222 308218 270986 308454
rect 271222 308218 306986 308454
rect 307222 308218 342986 308454
rect 343222 308218 378986 308454
rect 379222 308218 414986 308454
rect 415222 308218 450986 308454
rect 451222 308218 486986 308454
rect 487222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586442 308454
rect 586678 308218 586860 308454
rect -2936 308134 586860 308218
rect -2936 307898 -2754 308134
rect -2518 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 90986 308134
rect 91222 307898 126986 308134
rect 127222 307898 162986 308134
rect 163222 307898 198986 308134
rect 199222 307898 234986 308134
rect 235222 307898 270986 308134
rect 271222 307898 306986 308134
rect 307222 307898 342986 308134
rect 343222 307898 378986 308134
rect 379222 307898 414986 308134
rect 415222 307898 450986 308134
rect 451222 307898 486986 308134
rect 487222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586442 308134
rect 586678 307898 586860 308134
rect -2936 307876 586860 307898
rect -2936 307874 -2336 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 90804 307874 91404 307876
rect 126804 307874 127404 307876
rect 162804 307874 163404 307876
rect 198804 307874 199404 307876
rect 234804 307874 235404 307876
rect 270804 307874 271404 307876
rect 306804 307874 307404 307876
rect 342804 307874 343404 307876
rect 378804 307874 379404 307876
rect 414804 307874 415404 307876
rect 450804 307874 451404 307876
rect 486804 307874 487404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586260 307874 586860 307876
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 108804 290476 109404 290478
rect 144804 290476 145404 290478
rect 180804 290476 181404 290478
rect 216804 290476 217404 290478
rect 252804 290476 253404 290478
rect 288804 290476 289404 290478
rect 324804 290476 325404 290478
rect 360804 290476 361404 290478
rect 396804 290476 397404 290478
rect 432804 290476 433404 290478
rect 468804 290476 469404 290478
rect 504804 290476 505404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2936 290454 586860 290476
rect -2936 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 108986 290454
rect 109222 290218 144986 290454
rect 145222 290218 180986 290454
rect 181222 290218 216986 290454
rect 217222 290218 252986 290454
rect 253222 290218 288986 290454
rect 289222 290218 324986 290454
rect 325222 290218 360986 290454
rect 361222 290218 396986 290454
rect 397222 290218 432986 290454
rect 433222 290218 468986 290454
rect 469222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586860 290454
rect -2936 290134 586860 290218
rect -2936 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 108986 290134
rect 109222 289898 144986 290134
rect 145222 289898 180986 290134
rect 181222 289898 216986 290134
rect 217222 289898 252986 290134
rect 253222 289898 288986 290134
rect 289222 289898 324986 290134
rect 325222 289898 360986 290134
rect 361222 289898 396986 290134
rect 397222 289898 432986 290134
rect 433222 289898 468986 290134
rect 469222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586860 290134
rect -2936 289876 586860 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 108804 289874 109404 289876
rect 144804 289874 145404 289876
rect 180804 289874 181404 289876
rect 216804 289874 217404 289876
rect 252804 289874 253404 289876
rect 288804 289874 289404 289876
rect 324804 289874 325404 289876
rect 360804 289874 361404 289876
rect 396804 289874 397404 289876
rect 432804 289874 433404 289876
rect 468804 289874 469404 289876
rect 504804 289874 505404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -2936 272476 -2336 272478
rect 18804 272476 19404 272478
rect 270804 272476 271404 272478
rect 306804 272476 307404 272478
rect 586260 272476 586860 272478
rect -2936 272454 586860 272476
rect -2936 272218 -2754 272454
rect -2518 272218 18986 272454
rect 19222 272218 270986 272454
rect 271222 272218 306986 272454
rect 307222 272218 586442 272454
rect 586678 272218 586860 272454
rect -2936 272134 586860 272218
rect -2936 271898 -2754 272134
rect -2518 271898 18986 272134
rect 19222 271898 270986 272134
rect 271222 271898 306986 272134
rect 307222 271898 586442 272134
rect 586678 271898 586860 272134
rect -2936 271876 586860 271898
rect -2936 271874 -2336 271876
rect 18804 271874 19404 271876
rect 270804 271874 271404 271876
rect 306804 271874 307404 271876
rect 586260 271874 586860 271876
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 47088 254476 47408 254478
rect 77808 254476 78128 254478
rect 108528 254476 108848 254478
rect 139248 254476 139568 254478
rect 169968 254476 170288 254478
rect 200688 254476 201008 254478
rect 231408 254476 231728 254478
rect 262128 254476 262448 254478
rect 288804 254476 289404 254478
rect 339216 254476 339536 254478
rect 369936 254476 370256 254478
rect 400656 254476 400976 254478
rect 431376 254476 431696 254478
rect 462096 254476 462416 254478
rect 492816 254476 493136 254478
rect 523536 254476 523856 254478
rect 554256 254476 554576 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2936 254454 586860 254476
rect -2936 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 47130 254454
rect 47366 254218 77850 254454
rect 78086 254218 108570 254454
rect 108806 254218 139290 254454
rect 139526 254218 170010 254454
rect 170246 254218 200730 254454
rect 200966 254218 231450 254454
rect 231686 254218 262170 254454
rect 262406 254218 288986 254454
rect 289222 254218 339258 254454
rect 339494 254218 369978 254454
rect 370214 254218 400698 254454
rect 400934 254218 431418 254454
rect 431654 254218 462138 254454
rect 462374 254218 492858 254454
rect 493094 254218 523578 254454
rect 523814 254218 554298 254454
rect 554534 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586860 254454
rect -2936 254134 586860 254218
rect -2936 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 47130 254134
rect 47366 253898 77850 254134
rect 78086 253898 108570 254134
rect 108806 253898 139290 254134
rect 139526 253898 170010 254134
rect 170246 253898 200730 254134
rect 200966 253898 231450 254134
rect 231686 253898 262170 254134
rect 262406 253898 288986 254134
rect 289222 253898 339258 254134
rect 339494 253898 369978 254134
rect 370214 253898 400698 254134
rect 400934 253898 431418 254134
rect 431654 253898 462138 254134
rect 462374 253898 492858 254134
rect 493094 253898 523578 254134
rect 523814 253898 554298 254134
rect 554534 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586860 254134
rect -2936 253876 586860 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 47088 253874 47408 253876
rect 77808 253874 78128 253876
rect 108528 253874 108848 253876
rect 139248 253874 139568 253876
rect 169968 253874 170288 253876
rect 200688 253874 201008 253876
rect 231408 253874 231728 253876
rect 262128 253874 262448 253876
rect 288804 253874 289404 253876
rect 339216 253874 339536 253876
rect 369936 253874 370256 253876
rect 400656 253874 400976 253876
rect 431376 253874 431696 253876
rect 462096 253874 462416 253876
rect 492816 253874 493136 253876
rect 523536 253874 523856 253876
rect 554256 253874 554576 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -2936 236476 -2336 236478
rect 18804 236476 19404 236478
rect 31728 236476 32048 236478
rect 62448 236476 62768 236478
rect 93168 236476 93488 236478
rect 123888 236476 124208 236478
rect 154608 236476 154928 236478
rect 185328 236476 185648 236478
rect 216048 236476 216368 236478
rect 246768 236476 247088 236478
rect 270804 236476 271404 236478
rect 306804 236476 307404 236478
rect 323856 236476 324176 236478
rect 354576 236476 354896 236478
rect 385296 236476 385616 236478
rect 416016 236476 416336 236478
rect 446736 236476 447056 236478
rect 477456 236476 477776 236478
rect 508176 236476 508496 236478
rect 538896 236476 539216 236478
rect 586260 236476 586860 236478
rect -2936 236454 586860 236476
rect -2936 236218 -2754 236454
rect -2518 236218 18986 236454
rect 19222 236218 31770 236454
rect 32006 236218 62490 236454
rect 62726 236218 93210 236454
rect 93446 236218 123930 236454
rect 124166 236218 154650 236454
rect 154886 236218 185370 236454
rect 185606 236218 216090 236454
rect 216326 236218 246810 236454
rect 247046 236218 270986 236454
rect 271222 236218 306986 236454
rect 307222 236218 323898 236454
rect 324134 236218 354618 236454
rect 354854 236218 385338 236454
rect 385574 236218 416058 236454
rect 416294 236218 446778 236454
rect 447014 236218 477498 236454
rect 477734 236218 508218 236454
rect 508454 236218 538938 236454
rect 539174 236218 586442 236454
rect 586678 236218 586860 236454
rect -2936 236134 586860 236218
rect -2936 235898 -2754 236134
rect -2518 235898 18986 236134
rect 19222 235898 31770 236134
rect 32006 235898 62490 236134
rect 62726 235898 93210 236134
rect 93446 235898 123930 236134
rect 124166 235898 154650 236134
rect 154886 235898 185370 236134
rect 185606 235898 216090 236134
rect 216326 235898 246810 236134
rect 247046 235898 270986 236134
rect 271222 235898 306986 236134
rect 307222 235898 323898 236134
rect 324134 235898 354618 236134
rect 354854 235898 385338 236134
rect 385574 235898 416058 236134
rect 416294 235898 446778 236134
rect 447014 235898 477498 236134
rect 477734 235898 508218 236134
rect 508454 235898 538938 236134
rect 539174 235898 586442 236134
rect 586678 235898 586860 236134
rect -2936 235876 586860 235898
rect -2936 235874 -2336 235876
rect 18804 235874 19404 235876
rect 31728 235874 32048 235876
rect 62448 235874 62768 235876
rect 93168 235874 93488 235876
rect 123888 235874 124208 235876
rect 154608 235874 154928 235876
rect 185328 235874 185648 235876
rect 216048 235874 216368 235876
rect 246768 235874 247088 235876
rect 270804 235874 271404 235876
rect 306804 235874 307404 235876
rect 323856 235874 324176 235876
rect 354576 235874 354896 235876
rect 385296 235874 385616 235876
rect 416016 235874 416336 235876
rect 446736 235874 447056 235876
rect 477456 235874 477776 235876
rect 508176 235874 508496 235876
rect 538896 235874 539216 235876
rect 586260 235874 586860 235876
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 47088 218476 47408 218478
rect 77808 218476 78128 218478
rect 108528 218476 108848 218478
rect 139248 218476 139568 218478
rect 169968 218476 170288 218478
rect 200688 218476 201008 218478
rect 231408 218476 231728 218478
rect 262128 218476 262448 218478
rect 288804 218476 289404 218478
rect 339216 218476 339536 218478
rect 369936 218476 370256 218478
rect 400656 218476 400976 218478
rect 431376 218476 431696 218478
rect 462096 218476 462416 218478
rect 492816 218476 493136 218478
rect 523536 218476 523856 218478
rect 554256 218476 554576 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2936 218454 586860 218476
rect -2936 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 47130 218454
rect 47366 218218 77850 218454
rect 78086 218218 108570 218454
rect 108806 218218 139290 218454
rect 139526 218218 170010 218454
rect 170246 218218 200730 218454
rect 200966 218218 231450 218454
rect 231686 218218 262170 218454
rect 262406 218218 288986 218454
rect 289222 218218 339258 218454
rect 339494 218218 369978 218454
rect 370214 218218 400698 218454
rect 400934 218218 431418 218454
rect 431654 218218 462138 218454
rect 462374 218218 492858 218454
rect 493094 218218 523578 218454
rect 523814 218218 554298 218454
rect 554534 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586860 218454
rect -2936 218134 586860 218218
rect -2936 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 47130 218134
rect 47366 217898 77850 218134
rect 78086 217898 108570 218134
rect 108806 217898 139290 218134
rect 139526 217898 170010 218134
rect 170246 217898 200730 218134
rect 200966 217898 231450 218134
rect 231686 217898 262170 218134
rect 262406 217898 288986 218134
rect 289222 217898 339258 218134
rect 339494 217898 369978 218134
rect 370214 217898 400698 218134
rect 400934 217898 431418 218134
rect 431654 217898 462138 218134
rect 462374 217898 492858 218134
rect 493094 217898 523578 218134
rect 523814 217898 554298 218134
rect 554534 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586860 218134
rect -2936 217876 586860 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 47088 217874 47408 217876
rect 77808 217874 78128 217876
rect 108528 217874 108848 217876
rect 139248 217874 139568 217876
rect 169968 217874 170288 217876
rect 200688 217874 201008 217876
rect 231408 217874 231728 217876
rect 262128 217874 262448 217876
rect 288804 217874 289404 217876
rect 339216 217874 339536 217876
rect 369936 217874 370256 217876
rect 400656 217874 400976 217876
rect 431376 217874 431696 217876
rect 462096 217874 462416 217876
rect 492816 217874 493136 217876
rect 523536 217874 523856 217876
rect 554256 217874 554576 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -2936 200476 -2336 200478
rect 18804 200476 19404 200478
rect 31728 200476 32048 200478
rect 62448 200476 62768 200478
rect 93168 200476 93488 200478
rect 123888 200476 124208 200478
rect 154608 200476 154928 200478
rect 185328 200476 185648 200478
rect 216048 200476 216368 200478
rect 246768 200476 247088 200478
rect 270804 200476 271404 200478
rect 306804 200476 307404 200478
rect 323856 200476 324176 200478
rect 354576 200476 354896 200478
rect 385296 200476 385616 200478
rect 416016 200476 416336 200478
rect 446736 200476 447056 200478
rect 477456 200476 477776 200478
rect 508176 200476 508496 200478
rect 538896 200476 539216 200478
rect 586260 200476 586860 200478
rect -2936 200454 586860 200476
rect -2936 200218 -2754 200454
rect -2518 200218 18986 200454
rect 19222 200218 31770 200454
rect 32006 200218 62490 200454
rect 62726 200218 93210 200454
rect 93446 200218 123930 200454
rect 124166 200218 154650 200454
rect 154886 200218 185370 200454
rect 185606 200218 216090 200454
rect 216326 200218 246810 200454
rect 247046 200218 270986 200454
rect 271222 200218 306986 200454
rect 307222 200218 323898 200454
rect 324134 200218 354618 200454
rect 354854 200218 385338 200454
rect 385574 200218 416058 200454
rect 416294 200218 446778 200454
rect 447014 200218 477498 200454
rect 477734 200218 508218 200454
rect 508454 200218 538938 200454
rect 539174 200218 586442 200454
rect 586678 200218 586860 200454
rect -2936 200134 586860 200218
rect -2936 199898 -2754 200134
rect -2518 199898 18986 200134
rect 19222 199898 31770 200134
rect 32006 199898 62490 200134
rect 62726 199898 93210 200134
rect 93446 199898 123930 200134
rect 124166 199898 154650 200134
rect 154886 199898 185370 200134
rect 185606 199898 216090 200134
rect 216326 199898 246810 200134
rect 247046 199898 270986 200134
rect 271222 199898 306986 200134
rect 307222 199898 323898 200134
rect 324134 199898 354618 200134
rect 354854 199898 385338 200134
rect 385574 199898 416058 200134
rect 416294 199898 446778 200134
rect 447014 199898 477498 200134
rect 477734 199898 508218 200134
rect 508454 199898 538938 200134
rect 539174 199898 586442 200134
rect 586678 199898 586860 200134
rect -2936 199876 586860 199898
rect -2936 199874 -2336 199876
rect 18804 199874 19404 199876
rect 31728 199874 32048 199876
rect 62448 199874 62768 199876
rect 93168 199874 93488 199876
rect 123888 199874 124208 199876
rect 154608 199874 154928 199876
rect 185328 199874 185648 199876
rect 216048 199874 216368 199876
rect 246768 199874 247088 199876
rect 270804 199874 271404 199876
rect 306804 199874 307404 199876
rect 323856 199874 324176 199876
rect 354576 199874 354896 199876
rect 385296 199874 385616 199876
rect 416016 199874 416336 199876
rect 446736 199874 447056 199876
rect 477456 199874 477776 199876
rect 508176 199874 508496 199876
rect 538896 199874 539216 199876
rect 586260 199874 586860 199876
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 47088 182476 47408 182478
rect 77808 182476 78128 182478
rect 108528 182476 108848 182478
rect 139248 182476 139568 182478
rect 169968 182476 170288 182478
rect 200688 182476 201008 182478
rect 231408 182476 231728 182478
rect 262128 182476 262448 182478
rect 288804 182476 289404 182478
rect 339216 182476 339536 182478
rect 369936 182476 370256 182478
rect 400656 182476 400976 182478
rect 431376 182476 431696 182478
rect 462096 182476 462416 182478
rect 492816 182476 493136 182478
rect 523536 182476 523856 182478
rect 554256 182476 554576 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2936 182454 586860 182476
rect -2936 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 47130 182454
rect 47366 182218 77850 182454
rect 78086 182218 108570 182454
rect 108806 182218 139290 182454
rect 139526 182218 170010 182454
rect 170246 182218 200730 182454
rect 200966 182218 231450 182454
rect 231686 182218 262170 182454
rect 262406 182218 288986 182454
rect 289222 182218 339258 182454
rect 339494 182218 369978 182454
rect 370214 182218 400698 182454
rect 400934 182218 431418 182454
rect 431654 182218 462138 182454
rect 462374 182218 492858 182454
rect 493094 182218 523578 182454
rect 523814 182218 554298 182454
rect 554534 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586860 182454
rect -2936 182134 586860 182218
rect -2936 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 47130 182134
rect 47366 181898 77850 182134
rect 78086 181898 108570 182134
rect 108806 181898 139290 182134
rect 139526 181898 170010 182134
rect 170246 181898 200730 182134
rect 200966 181898 231450 182134
rect 231686 181898 262170 182134
rect 262406 181898 288986 182134
rect 289222 181898 339258 182134
rect 339494 181898 369978 182134
rect 370214 181898 400698 182134
rect 400934 181898 431418 182134
rect 431654 181898 462138 182134
rect 462374 181898 492858 182134
rect 493094 181898 523578 182134
rect 523814 181898 554298 182134
rect 554534 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586860 182134
rect -2936 181876 586860 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 47088 181874 47408 181876
rect 77808 181874 78128 181876
rect 108528 181874 108848 181876
rect 139248 181874 139568 181876
rect 169968 181874 170288 181876
rect 200688 181874 201008 181876
rect 231408 181874 231728 181876
rect 262128 181874 262448 181876
rect 288804 181874 289404 181876
rect 339216 181874 339536 181876
rect 369936 181874 370256 181876
rect 400656 181874 400976 181876
rect 431376 181874 431696 181876
rect 462096 181874 462416 181876
rect 492816 181874 493136 181876
rect 523536 181874 523856 181876
rect 554256 181874 554576 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -2936 164476 -2336 164478
rect 18804 164476 19404 164478
rect 31728 164476 32048 164478
rect 62448 164476 62768 164478
rect 93168 164476 93488 164478
rect 123888 164476 124208 164478
rect 154608 164476 154928 164478
rect 185328 164476 185648 164478
rect 216048 164476 216368 164478
rect 246768 164476 247088 164478
rect 270804 164476 271404 164478
rect 306804 164476 307404 164478
rect 323856 164476 324176 164478
rect 354576 164476 354896 164478
rect 385296 164476 385616 164478
rect 416016 164476 416336 164478
rect 446736 164476 447056 164478
rect 477456 164476 477776 164478
rect 508176 164476 508496 164478
rect 538896 164476 539216 164478
rect 586260 164476 586860 164478
rect -2936 164454 586860 164476
rect -2936 164218 -2754 164454
rect -2518 164218 18986 164454
rect 19222 164218 31770 164454
rect 32006 164218 62490 164454
rect 62726 164218 93210 164454
rect 93446 164218 123930 164454
rect 124166 164218 154650 164454
rect 154886 164218 185370 164454
rect 185606 164218 216090 164454
rect 216326 164218 246810 164454
rect 247046 164218 270986 164454
rect 271222 164218 306986 164454
rect 307222 164218 323898 164454
rect 324134 164218 354618 164454
rect 354854 164218 385338 164454
rect 385574 164218 416058 164454
rect 416294 164218 446778 164454
rect 447014 164218 477498 164454
rect 477734 164218 508218 164454
rect 508454 164218 538938 164454
rect 539174 164218 586442 164454
rect 586678 164218 586860 164454
rect -2936 164134 586860 164218
rect -2936 163898 -2754 164134
rect -2518 163898 18986 164134
rect 19222 163898 31770 164134
rect 32006 163898 62490 164134
rect 62726 163898 93210 164134
rect 93446 163898 123930 164134
rect 124166 163898 154650 164134
rect 154886 163898 185370 164134
rect 185606 163898 216090 164134
rect 216326 163898 246810 164134
rect 247046 163898 270986 164134
rect 271222 163898 306986 164134
rect 307222 163898 323898 164134
rect 324134 163898 354618 164134
rect 354854 163898 385338 164134
rect 385574 163898 416058 164134
rect 416294 163898 446778 164134
rect 447014 163898 477498 164134
rect 477734 163898 508218 164134
rect 508454 163898 538938 164134
rect 539174 163898 586442 164134
rect 586678 163898 586860 164134
rect -2936 163876 586860 163898
rect -2936 163874 -2336 163876
rect 18804 163874 19404 163876
rect 31728 163874 32048 163876
rect 62448 163874 62768 163876
rect 93168 163874 93488 163876
rect 123888 163874 124208 163876
rect 154608 163874 154928 163876
rect 185328 163874 185648 163876
rect 216048 163874 216368 163876
rect 246768 163874 247088 163876
rect 270804 163874 271404 163876
rect 306804 163874 307404 163876
rect 323856 163874 324176 163876
rect 354576 163874 354896 163876
rect 385296 163874 385616 163876
rect 416016 163874 416336 163876
rect 446736 163874 447056 163876
rect 477456 163874 477776 163876
rect 508176 163874 508496 163876
rect 538896 163874 539216 163876
rect 586260 163874 586860 163876
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 47088 146476 47408 146478
rect 77808 146476 78128 146478
rect 108528 146476 108848 146478
rect 139248 146476 139568 146478
rect 169968 146476 170288 146478
rect 200688 146476 201008 146478
rect 231408 146476 231728 146478
rect 262128 146476 262448 146478
rect 288804 146476 289404 146478
rect 339216 146476 339536 146478
rect 369936 146476 370256 146478
rect 400656 146476 400976 146478
rect 431376 146476 431696 146478
rect 462096 146476 462416 146478
rect 492816 146476 493136 146478
rect 523536 146476 523856 146478
rect 554256 146476 554576 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2936 146454 586860 146476
rect -2936 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 47130 146454
rect 47366 146218 77850 146454
rect 78086 146218 108570 146454
rect 108806 146218 139290 146454
rect 139526 146218 170010 146454
rect 170246 146218 200730 146454
rect 200966 146218 231450 146454
rect 231686 146218 262170 146454
rect 262406 146218 288986 146454
rect 289222 146218 339258 146454
rect 339494 146218 369978 146454
rect 370214 146218 400698 146454
rect 400934 146218 431418 146454
rect 431654 146218 462138 146454
rect 462374 146218 492858 146454
rect 493094 146218 523578 146454
rect 523814 146218 554298 146454
rect 554534 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586860 146454
rect -2936 146134 586860 146218
rect -2936 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 47130 146134
rect 47366 145898 77850 146134
rect 78086 145898 108570 146134
rect 108806 145898 139290 146134
rect 139526 145898 170010 146134
rect 170246 145898 200730 146134
rect 200966 145898 231450 146134
rect 231686 145898 262170 146134
rect 262406 145898 288986 146134
rect 289222 145898 339258 146134
rect 339494 145898 369978 146134
rect 370214 145898 400698 146134
rect 400934 145898 431418 146134
rect 431654 145898 462138 146134
rect 462374 145898 492858 146134
rect 493094 145898 523578 146134
rect 523814 145898 554298 146134
rect 554534 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586860 146134
rect -2936 145876 586860 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 47088 145874 47408 145876
rect 77808 145874 78128 145876
rect 108528 145874 108848 145876
rect 139248 145874 139568 145876
rect 169968 145874 170288 145876
rect 200688 145874 201008 145876
rect 231408 145874 231728 145876
rect 262128 145874 262448 145876
rect 288804 145874 289404 145876
rect 339216 145874 339536 145876
rect 369936 145874 370256 145876
rect 400656 145874 400976 145876
rect 431376 145874 431696 145876
rect 462096 145874 462416 145876
rect 492816 145874 493136 145876
rect 523536 145874 523856 145876
rect 554256 145874 554576 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -2936 128476 -2336 128478
rect 18804 128476 19404 128478
rect 31728 128476 32048 128478
rect 62448 128476 62768 128478
rect 93168 128476 93488 128478
rect 123888 128476 124208 128478
rect 154608 128476 154928 128478
rect 185328 128476 185648 128478
rect 216048 128476 216368 128478
rect 246768 128476 247088 128478
rect 270804 128476 271404 128478
rect 306804 128476 307404 128478
rect 323856 128476 324176 128478
rect 354576 128476 354896 128478
rect 385296 128476 385616 128478
rect 416016 128476 416336 128478
rect 446736 128476 447056 128478
rect 477456 128476 477776 128478
rect 508176 128476 508496 128478
rect 538896 128476 539216 128478
rect 586260 128476 586860 128478
rect -2936 128454 586860 128476
rect -2936 128218 -2754 128454
rect -2518 128218 18986 128454
rect 19222 128218 31770 128454
rect 32006 128218 62490 128454
rect 62726 128218 93210 128454
rect 93446 128218 123930 128454
rect 124166 128218 154650 128454
rect 154886 128218 185370 128454
rect 185606 128218 216090 128454
rect 216326 128218 246810 128454
rect 247046 128218 270986 128454
rect 271222 128218 306986 128454
rect 307222 128218 323898 128454
rect 324134 128218 354618 128454
rect 354854 128218 385338 128454
rect 385574 128218 416058 128454
rect 416294 128218 446778 128454
rect 447014 128218 477498 128454
rect 477734 128218 508218 128454
rect 508454 128218 538938 128454
rect 539174 128218 586442 128454
rect 586678 128218 586860 128454
rect -2936 128134 586860 128218
rect -2936 127898 -2754 128134
rect -2518 127898 18986 128134
rect 19222 127898 31770 128134
rect 32006 127898 62490 128134
rect 62726 127898 93210 128134
rect 93446 127898 123930 128134
rect 124166 127898 154650 128134
rect 154886 127898 185370 128134
rect 185606 127898 216090 128134
rect 216326 127898 246810 128134
rect 247046 127898 270986 128134
rect 271222 127898 306986 128134
rect 307222 127898 323898 128134
rect 324134 127898 354618 128134
rect 354854 127898 385338 128134
rect 385574 127898 416058 128134
rect 416294 127898 446778 128134
rect 447014 127898 477498 128134
rect 477734 127898 508218 128134
rect 508454 127898 538938 128134
rect 539174 127898 586442 128134
rect 586678 127898 586860 128134
rect -2936 127876 586860 127898
rect -2936 127874 -2336 127876
rect 18804 127874 19404 127876
rect 31728 127874 32048 127876
rect 62448 127874 62768 127876
rect 93168 127874 93488 127876
rect 123888 127874 124208 127876
rect 154608 127874 154928 127876
rect 185328 127874 185648 127876
rect 216048 127874 216368 127876
rect 246768 127874 247088 127876
rect 270804 127874 271404 127876
rect 306804 127874 307404 127876
rect 323856 127874 324176 127876
rect 354576 127874 354896 127876
rect 385296 127874 385616 127876
rect 416016 127874 416336 127876
rect 446736 127874 447056 127876
rect 477456 127874 477776 127876
rect 508176 127874 508496 127876
rect 538896 127874 539216 127876
rect 586260 127874 586860 127876
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 47088 110476 47408 110478
rect 77808 110476 78128 110478
rect 108528 110476 108848 110478
rect 139248 110476 139568 110478
rect 169968 110476 170288 110478
rect 200688 110476 201008 110478
rect 231408 110476 231728 110478
rect 262128 110476 262448 110478
rect 288804 110476 289404 110478
rect 339216 110476 339536 110478
rect 369936 110476 370256 110478
rect 400656 110476 400976 110478
rect 431376 110476 431696 110478
rect 462096 110476 462416 110478
rect 492816 110476 493136 110478
rect 523536 110476 523856 110478
rect 554256 110476 554576 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2936 110454 586860 110476
rect -2936 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 47130 110454
rect 47366 110218 77850 110454
rect 78086 110218 108570 110454
rect 108806 110218 139290 110454
rect 139526 110218 170010 110454
rect 170246 110218 200730 110454
rect 200966 110218 231450 110454
rect 231686 110218 262170 110454
rect 262406 110218 288986 110454
rect 289222 110218 339258 110454
rect 339494 110218 369978 110454
rect 370214 110218 400698 110454
rect 400934 110218 431418 110454
rect 431654 110218 462138 110454
rect 462374 110218 492858 110454
rect 493094 110218 523578 110454
rect 523814 110218 554298 110454
rect 554534 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586860 110454
rect -2936 110134 586860 110218
rect -2936 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 47130 110134
rect 47366 109898 77850 110134
rect 78086 109898 108570 110134
rect 108806 109898 139290 110134
rect 139526 109898 170010 110134
rect 170246 109898 200730 110134
rect 200966 109898 231450 110134
rect 231686 109898 262170 110134
rect 262406 109898 288986 110134
rect 289222 109898 339258 110134
rect 339494 109898 369978 110134
rect 370214 109898 400698 110134
rect 400934 109898 431418 110134
rect 431654 109898 462138 110134
rect 462374 109898 492858 110134
rect 493094 109898 523578 110134
rect 523814 109898 554298 110134
rect 554534 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586860 110134
rect -2936 109876 586860 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 47088 109874 47408 109876
rect 77808 109874 78128 109876
rect 108528 109874 108848 109876
rect 139248 109874 139568 109876
rect 169968 109874 170288 109876
rect 200688 109874 201008 109876
rect 231408 109874 231728 109876
rect 262128 109874 262448 109876
rect 288804 109874 289404 109876
rect 339216 109874 339536 109876
rect 369936 109874 370256 109876
rect 400656 109874 400976 109876
rect 431376 109874 431696 109876
rect 462096 109874 462416 109876
rect 492816 109874 493136 109876
rect 523536 109874 523856 109876
rect 554256 109874 554576 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -2936 92476 -2336 92478
rect 18804 92476 19404 92478
rect 31728 92476 32048 92478
rect 62448 92476 62768 92478
rect 93168 92476 93488 92478
rect 123888 92476 124208 92478
rect 154608 92476 154928 92478
rect 185328 92476 185648 92478
rect 216048 92476 216368 92478
rect 246768 92476 247088 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 323856 92476 324176 92478
rect 354576 92476 354896 92478
rect 385296 92476 385616 92478
rect 416016 92476 416336 92478
rect 446736 92476 447056 92478
rect 477456 92476 477776 92478
rect 508176 92476 508496 92478
rect 538896 92476 539216 92478
rect 586260 92476 586860 92478
rect -2936 92454 586860 92476
rect -2936 92218 -2754 92454
rect -2518 92218 18986 92454
rect 19222 92218 31770 92454
rect 32006 92218 62490 92454
rect 62726 92218 93210 92454
rect 93446 92218 123930 92454
rect 124166 92218 154650 92454
rect 154886 92218 185370 92454
rect 185606 92218 216090 92454
rect 216326 92218 246810 92454
rect 247046 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 323898 92454
rect 324134 92218 354618 92454
rect 354854 92218 385338 92454
rect 385574 92218 416058 92454
rect 416294 92218 446778 92454
rect 447014 92218 477498 92454
rect 477734 92218 508218 92454
rect 508454 92218 538938 92454
rect 539174 92218 586442 92454
rect 586678 92218 586860 92454
rect -2936 92134 586860 92218
rect -2936 91898 -2754 92134
rect -2518 91898 18986 92134
rect 19222 91898 31770 92134
rect 32006 91898 62490 92134
rect 62726 91898 93210 92134
rect 93446 91898 123930 92134
rect 124166 91898 154650 92134
rect 154886 91898 185370 92134
rect 185606 91898 216090 92134
rect 216326 91898 246810 92134
rect 247046 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 323898 92134
rect 324134 91898 354618 92134
rect 354854 91898 385338 92134
rect 385574 91898 416058 92134
rect 416294 91898 446778 92134
rect 447014 91898 477498 92134
rect 477734 91898 508218 92134
rect 508454 91898 538938 92134
rect 539174 91898 586442 92134
rect 586678 91898 586860 92134
rect -2936 91876 586860 91898
rect -2936 91874 -2336 91876
rect 18804 91874 19404 91876
rect 31728 91874 32048 91876
rect 62448 91874 62768 91876
rect 93168 91874 93488 91876
rect 123888 91874 124208 91876
rect 154608 91874 154928 91876
rect 185328 91874 185648 91876
rect 216048 91874 216368 91876
rect 246768 91874 247088 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 323856 91874 324176 91876
rect 354576 91874 354896 91876
rect 385296 91874 385616 91876
rect 416016 91874 416336 91876
rect 446736 91874 447056 91876
rect 477456 91874 477776 91876
rect 508176 91874 508496 91876
rect 538896 91874 539216 91876
rect 586260 91874 586860 91876
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 288804 74476 289404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2936 74454 586860 74476
rect -2936 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 288986 74454
rect 289222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586860 74454
rect -2936 74134 586860 74218
rect -2936 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 288986 74134
rect 289222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586860 74134
rect -2936 73876 586860 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 288804 73874 289404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -2936 56476 -2336 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586260 56476 586860 56478
rect -2936 56454 586860 56476
rect -2936 56218 -2754 56454
rect -2518 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586442 56454
rect 586678 56218 586860 56454
rect -2936 56134 586860 56218
rect -2936 55898 -2754 56134
rect -2518 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586442 56134
rect 586678 55898 586860 56134
rect -2936 55876 586860 55898
rect -2936 55874 -2336 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586260 55874 586860 55876
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2936 38454 586860 38476
rect -2936 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586860 38454
rect -2936 38134 586860 38218
rect -2936 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586860 38134
rect -2936 37876 586860 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -2936 20476 -2336 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586260 20476 586860 20478
rect -2936 20454 586860 20476
rect -2936 20218 -2754 20454
rect -2518 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586442 20454
rect 586678 20218 586860 20454
rect -2936 20134 586860 20218
rect -2936 19898 -2754 20134
rect -2518 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586442 20134
rect 586678 19898 586860 20134
rect -2936 19876 586860 19898
rect -2936 19874 -2336 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586260 19874 586860 19876
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2936 2454 586860 2476
rect -2936 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586860 2454
rect -2936 2134 586860 2218
rect -2936 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586860 2134
rect -2936 1876 586860 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 18804 -1264 19404 -1262
rect 54804 -1264 55404 -1262
rect 90804 -1264 91404 -1262
rect 126804 -1264 127404 -1262
rect 162804 -1264 163404 -1262
rect 198804 -1264 199404 -1262
rect 234804 -1264 235404 -1262
rect 270804 -1264 271404 -1262
rect 306804 -1264 307404 -1262
rect 342804 -1264 343404 -1262
rect 378804 -1264 379404 -1262
rect 414804 -1264 415404 -1262
rect 450804 -1264 451404 -1262
rect 486804 -1264 487404 -1262
rect 522804 -1264 523404 -1262
rect 558804 -1264 559404 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1286 586860 -1264
rect -2936 -1522 -2754 -1286
rect -2518 -1522 18986 -1286
rect 19222 -1522 54986 -1286
rect 55222 -1522 90986 -1286
rect 91222 -1522 126986 -1286
rect 127222 -1522 162986 -1286
rect 163222 -1522 198986 -1286
rect 199222 -1522 234986 -1286
rect 235222 -1522 270986 -1286
rect 271222 -1522 306986 -1286
rect 307222 -1522 342986 -1286
rect 343222 -1522 378986 -1286
rect 379222 -1522 414986 -1286
rect 415222 -1522 450986 -1286
rect 451222 -1522 486986 -1286
rect 487222 -1522 522986 -1286
rect 523222 -1522 558986 -1286
rect 559222 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect -2936 -1606 586860 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 18986 -1606
rect 19222 -1842 54986 -1606
rect 55222 -1842 90986 -1606
rect 91222 -1842 126986 -1606
rect 127222 -1842 162986 -1606
rect 163222 -1842 198986 -1606
rect 199222 -1842 234986 -1606
rect 235222 -1842 270986 -1606
rect 271222 -1842 306986 -1606
rect 307222 -1842 342986 -1606
rect 343222 -1842 378986 -1606
rect 379222 -1842 414986 -1606
rect 415222 -1842 450986 -1606
rect 451222 -1842 486986 -1606
rect 487222 -1842 522986 -1606
rect 523222 -1842 558986 -1606
rect 559222 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect -2936 -1864 586860 -1842
rect -2936 -1866 -2336 -1864
rect 18804 -1866 19404 -1864
rect 54804 -1866 55404 -1864
rect 90804 -1866 91404 -1864
rect 126804 -1866 127404 -1864
rect 162804 -1866 163404 -1864
rect 198804 -1866 199404 -1864
rect 234804 -1866 235404 -1864
rect 270804 -1866 271404 -1864
rect 306804 -1866 307404 -1864
rect 342804 -1866 343404 -1864
rect 378804 -1866 379404 -1864
rect 414804 -1866 415404 -1864
rect 450804 -1866 451404 -1864
rect 486804 -1866 487404 -1864
rect 522804 -1866 523404 -1864
rect 558804 -1866 559404 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2226 587800 -2204
rect -3876 -2462 -3694 -2226
rect -3458 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect -3876 -2546 587800 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect -3876 -2804 587800 -2782
rect -3876 -2806 -3276 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3166 588740 -3144
rect -4816 -3402 -4634 -3166
rect -4398 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect -4816 -3486 588740 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect -4816 -3744 588740 -3722
rect -4816 -3746 -4216 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4106 589680 -4084
rect -5756 -4342 -5574 -4106
rect -5338 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect -5756 -4426 589680 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect -5756 -4684 589680 -4662
rect -5756 -4686 -5156 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5046 590620 -5024
rect -6696 -5282 -6514 -5046
rect -6278 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect -6696 -5366 590620 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect -6696 -5624 590620 -5602
rect -6696 -5626 -6096 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 590960 -5964 591560 -5962
rect -7636 -5986 591560 -5964
rect -7636 -6222 -7454 -5986
rect -7218 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect -7636 -6306 591560 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect -7636 -6564 591560 -6542
rect -7636 -6566 -7036 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 591900 -6904 592500 -6902
rect -8576 -6926 592500 -6904
rect -8576 -7162 -8394 -6926
rect -8158 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect -8576 -7246 592500 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect -8576 -7504 592500 -7482
rect -8576 -7506 -7976 -7504
rect 591900 -7506 592500 -7504
use decred_hash_macro  decred_hash_block3
timestamp 1608259780
transform -1 0 558784 0 -1 583916
box 0 0 240000 200000
use decred_hash_macro  decred_hash_block2
timestamp 1608259780
transform -1 0 266656 0 -1 583916
box 0 0 240000 200000
use decred_hash_macro  decred_hash_block1
timestamp 1608259780
transform -1 0 558784 0 -1 273600
box 0 0 240000 200000
use decred_hash_macro  decred_hash_block0
timestamp 1608259780
transform -1 0 266656 0 -1 273600
box 0 0 240000 200000
use decred_controller  decred_controller_block
timestamp 1608259780
transform -1 0 312000 0 -1 355560
box 0 0 40000 40000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew signal bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew signal bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew signal bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew signal input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew signal input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew signal input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew signal input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew signal input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew signal input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew signal input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew signal input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew signal input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew signal input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew signal input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew signal input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew signal input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew signal input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew signal input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew signal input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew signal input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew signal input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew signal input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew signal input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew signal input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew signal input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew signal input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew signal input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew signal input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew signal input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew signal input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew signal input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew signal input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew signal tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 70 nsew signal tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 71 nsew signal tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 72 nsew signal tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 73 nsew signal tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 74 nsew signal tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 75 nsew signal tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 76 nsew signal tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 77 nsew signal tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 78 nsew signal tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 79 nsew signal tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 80 nsew signal tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 81 nsew signal tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 82 nsew signal tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 83 nsew signal tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 84 nsew signal tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 85 nsew signal tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 86 nsew signal tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 87 nsew signal tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 88 nsew signal tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 89 nsew signal tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 90 nsew signal tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 91 nsew signal tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 92 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 93 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 94 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 95 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 96 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 97 nsew signal tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 98 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 99 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 100 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 101 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 102 nsew signal tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 103 nsew signal tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 104 nsew signal tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 105 nsew signal tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 106 nsew signal tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 107 nsew signal tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 108 nsew signal tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 109 nsew signal tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 110 nsew signal tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 111 nsew signal tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 112 nsew signal tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 113 nsew signal tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 114 nsew signal tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 115 nsew signal tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 116 nsew signal tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 117 nsew signal tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 118 nsew signal tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 119 nsew signal tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 120 nsew signal tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 121 nsew signal tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 122 nsew signal tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 123 nsew signal tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 124 nsew signal tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 125 nsew signal input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 126 nsew signal input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 127 nsew signal input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 128 nsew signal input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 129 nsew signal input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 130 nsew signal input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 131 nsew signal input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 132 nsew signal input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 133 nsew signal input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 134 nsew signal input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 135 nsew signal input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 136 nsew signal input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 137 nsew signal input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 138 nsew signal input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 139 nsew signal input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 140 nsew signal input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 141 nsew signal input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 142 nsew signal input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 143 nsew signal input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 144 nsew signal input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 145 nsew signal input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 146 nsew signal input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 147 nsew signal input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 148 nsew signal input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 149 nsew signal input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 150 nsew signal input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 151 nsew signal input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 152 nsew signal input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 153 nsew signal input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 154 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 155 nsew signal input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 156 nsew signal input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 157 nsew signal input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 158 nsew signal input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 159 nsew signal input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 160 nsew signal input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 161 nsew signal input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 162 nsew signal input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 163 nsew signal input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 164 nsew signal input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 165 nsew signal input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 166 nsew signal input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 167 nsew signal input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 168 nsew signal input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 169 nsew signal input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 170 nsew signal input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 171 nsew signal input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 172 nsew signal input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 173 nsew signal input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 174 nsew signal input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 175 nsew signal input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 176 nsew signal input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 177 nsew signal input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 178 nsew signal input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 179 nsew signal input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 180 nsew signal input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 181 nsew signal input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 182 nsew signal input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 183 nsew signal input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 184 nsew signal input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 185 nsew signal input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 186 nsew signal input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 187 nsew signal input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 188 nsew signal input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 189 nsew signal input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 190 nsew signal input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 191 nsew signal input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 192 nsew signal input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 193 nsew signal input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 194 nsew signal input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 195 nsew signal input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 196 nsew signal input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 197 nsew signal input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 198 nsew signal input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 199 nsew signal input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 200 nsew signal input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 201 nsew signal input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 202 nsew signal input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 203 nsew signal input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 204 nsew signal input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 205 nsew signal input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 206 nsew signal input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 207 nsew signal input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 208 nsew signal input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 209 nsew signal input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 210 nsew signal input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 211 nsew signal input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 212 nsew signal input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 213 nsew signal input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 214 nsew signal input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 215 nsew signal input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 216 nsew signal input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 217 nsew signal input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 218 nsew signal input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 219 nsew signal input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 220 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 221 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 222 nsew signal input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 223 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 224 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 225 nsew signal input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 226 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 227 nsew signal input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 228 nsew signal input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 229 nsew signal input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 230 nsew signal input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 231 nsew signal input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 232 nsew signal input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 233 nsew signal input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 234 nsew signal input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 235 nsew signal input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 236 nsew signal input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 237 nsew signal input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 238 nsew signal input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 239 nsew signal input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 240 nsew signal input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 241 nsew signal input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 242 nsew signal input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 243 nsew signal input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 244 nsew signal input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 245 nsew signal input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 246 nsew signal input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 247 nsew signal input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 248 nsew signal input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 249 nsew signal input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 250 nsew signal input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 251 nsew signal input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 252 nsew signal input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 253 nsew signal tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 254 nsew signal tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 255 nsew signal tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 256 nsew signal tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 257 nsew signal tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 258 nsew signal tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 259 nsew signal tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 260 nsew signal tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 261 nsew signal tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 262 nsew signal tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 263 nsew signal tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 264 nsew signal tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 265 nsew signal tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 266 nsew signal tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 267 nsew signal tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 268 nsew signal tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 269 nsew signal tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 270 nsew signal tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 271 nsew signal tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 272 nsew signal tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 273 nsew signal tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 274 nsew signal tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 275 nsew signal tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 276 nsew signal tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 277 nsew signal tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 278 nsew signal tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 279 nsew signal tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 280 nsew signal tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 281 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 282 nsew signal tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 283 nsew signal tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 284 nsew signal tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 285 nsew signal tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 286 nsew signal tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 287 nsew signal tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 288 nsew signal tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 289 nsew signal tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 290 nsew signal tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 291 nsew signal tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 292 nsew signal tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 293 nsew signal tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 294 nsew signal tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 295 nsew signal tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 296 nsew signal tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 297 nsew signal tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 298 nsew signal tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 299 nsew signal tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 300 nsew signal tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 301 nsew signal tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 302 nsew signal tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 303 nsew signal tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 304 nsew signal tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 305 nsew signal tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 306 nsew signal tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 307 nsew signal tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 308 nsew signal tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 309 nsew signal tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 310 nsew signal tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 311 nsew signal tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 312 nsew signal tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 313 nsew signal tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 314 nsew signal tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 315 nsew signal tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 316 nsew signal tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 317 nsew signal tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 318 nsew signal tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 319 nsew signal tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 320 nsew signal tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 321 nsew signal tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 322 nsew signal tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 323 nsew signal tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 324 nsew signal tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 325 nsew signal tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 326 nsew signal tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 327 nsew signal tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 328 nsew signal tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 329 nsew signal tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 330 nsew signal tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 331 nsew signal tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 332 nsew signal tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 333 nsew signal tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 334 nsew signal tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 335 nsew signal tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 336 nsew signal tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 337 nsew signal tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 338 nsew signal tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 339 nsew signal tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 340 nsew signal tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 341 nsew signal tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 342 nsew signal tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 343 nsew signal tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 344 nsew signal tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 345 nsew signal tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 346 nsew signal tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 347 nsew signal tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 348 nsew signal tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 349 nsew signal tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 350 nsew signal tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 351 nsew signal tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 352 nsew signal tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 353 nsew signal tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 354 nsew signal tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 355 nsew signal tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 356 nsew signal tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 357 nsew signal tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 358 nsew signal tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 359 nsew signal tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 360 nsew signal tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 361 nsew signal tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 362 nsew signal tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 363 nsew signal tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 364 nsew signal tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 365 nsew signal tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 366 nsew signal tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 367 nsew signal tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 368 nsew signal tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 369 nsew signal tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 370 nsew signal tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 371 nsew signal tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 372 nsew signal tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 373 nsew signal tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 374 nsew signal tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 375 nsew signal tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 376 nsew signal tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 377 nsew signal tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 378 nsew signal tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 379 nsew signal tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 380 nsew signal tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 381 nsew signal input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 382 nsew signal input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 383 nsew signal input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 384 nsew signal input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 385 nsew signal input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 386 nsew signal input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 387 nsew signal input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 388 nsew signal input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 389 nsew signal input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 390 nsew signal input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 391 nsew signal input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 392 nsew signal input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 393 nsew signal input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 394 nsew signal input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 395 nsew signal input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 396 nsew signal input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 397 nsew signal input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 398 nsew signal input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 399 nsew signal input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 400 nsew signal input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 401 nsew signal input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 402 nsew signal input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 403 nsew signal input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 404 nsew signal input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 405 nsew signal input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 406 nsew signal input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 407 nsew signal input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 408 nsew signal input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 409 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 410 nsew signal input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 411 nsew signal input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 412 nsew signal input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 413 nsew signal input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 414 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 415 nsew signal input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 416 nsew signal input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 417 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 418 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 419 nsew signal input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 420 nsew signal input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 421 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 422 nsew signal input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 423 nsew signal input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 424 nsew signal input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 425 nsew signal input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 426 nsew signal input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 427 nsew signal input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 428 nsew signal input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 429 nsew signal input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 430 nsew signal input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 431 nsew signal input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 432 nsew signal input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 433 nsew signal input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 434 nsew signal input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 435 nsew signal input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 436 nsew signal input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 437 nsew signal input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 438 nsew signal input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 439 nsew signal input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 440 nsew signal input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 441 nsew signal input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 442 nsew signal input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 443 nsew signal input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 444 nsew signal input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 445 nsew signal input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 446 nsew signal input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 447 nsew signal input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 448 nsew signal input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 449 nsew signal input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 450 nsew signal input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 451 nsew signal input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 452 nsew signal input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 453 nsew signal input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 454 nsew signal input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 455 nsew signal input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 456 nsew signal input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 457 nsew signal input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 458 nsew signal input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 459 nsew signal input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 460 nsew signal input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 461 nsew signal input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 462 nsew signal input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 463 nsew signal input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 464 nsew signal input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 465 nsew signal input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 466 nsew signal input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 467 nsew signal input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 468 nsew signal input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 469 nsew signal input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 470 nsew signal input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 471 nsew signal input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 472 nsew signal input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 473 nsew signal input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 474 nsew signal input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 475 nsew signal input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 476 nsew signal input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 477 nsew signal input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 478 nsew signal input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 479 nsew signal input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 480 nsew signal input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 481 nsew signal input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 482 nsew signal input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 483 nsew signal input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 484 nsew signal input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 485 nsew signal input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 486 nsew signal input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 487 nsew signal input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 488 nsew signal input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 489 nsew signal input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 490 nsew signal input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 491 nsew signal input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 492 nsew signal input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 493 nsew signal input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 494 nsew signal input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 495 nsew signal input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 496 nsew signal input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 497 nsew signal input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 498 nsew signal input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 499 nsew signal input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 500 nsew signal input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 501 nsew signal input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 502 nsew signal input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 503 nsew signal input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 504 nsew signal input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 505 nsew signal input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 506 nsew signal input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 507 nsew signal input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 508 nsew signal input
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 509 nsew signal tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 510 nsew signal tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 511 nsew signal tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 512 nsew signal tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 513 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 514 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 515 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 516 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 517 nsew signal tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 518 nsew signal tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 519 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 520 nsew signal input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 521 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 522 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 523 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 524 nsew signal input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 525 nsew signal input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 526 nsew signal input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 527 nsew signal input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 528 nsew signal input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 529 nsew signal input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 530 nsew signal input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 531 nsew signal input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 532 nsew signal input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 533 nsew signal input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 534 nsew signal input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 535 nsew signal input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 536 nsew signal input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 537 nsew signal input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 538 nsew signal input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 539 nsew signal input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 540 nsew signal input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 541 nsew signal input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 542 nsew signal input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 543 nsew signal input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 544 nsew signal input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 545 nsew signal input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 546 nsew signal input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 547 nsew signal input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 548 nsew signal input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 549 nsew signal input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 550 nsew signal input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 551 nsew signal input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 552 nsew signal input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 553 nsew signal input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 554 nsew signal input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 555 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 556 nsew signal input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 557 nsew signal input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 558 nsew signal input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 559 nsew signal input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 560 nsew signal input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 561 nsew signal input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 562 nsew signal input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 563 nsew signal input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 564 nsew signal input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 565 nsew signal input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 566 nsew signal input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 567 nsew signal input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 568 nsew signal input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 569 nsew signal input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 570 nsew signal input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 571 nsew signal input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 572 nsew signal input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 573 nsew signal input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 574 nsew signal input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 575 nsew signal input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 576 nsew signal input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 577 nsew signal input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 578 nsew signal input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 579 nsew signal input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 580 nsew signal input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 581 nsew signal input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 582 nsew signal input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 583 nsew signal input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 584 nsew signal input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 585 nsew signal input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 586 nsew signal input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 587 nsew signal input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 588 nsew signal input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 589 nsew signal tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 590 nsew signal tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 591 nsew signal tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 592 nsew signal tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 593 nsew signal tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 594 nsew signal tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 595 nsew signal tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 596 nsew signal tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 597 nsew signal tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 598 nsew signal tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 599 nsew signal tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 600 nsew signal tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 601 nsew signal tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 602 nsew signal tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 603 nsew signal tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 604 nsew signal tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 605 nsew signal tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 606 nsew signal tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 607 nsew signal tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 608 nsew signal tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 609 nsew signal tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 610 nsew signal tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 611 nsew signal tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 612 nsew signal tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 613 nsew signal tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 614 nsew signal tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 615 nsew signal tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 616 nsew signal tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 617 nsew signal tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 618 nsew signal tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 619 nsew signal tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 620 nsew signal tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 621 nsew signal input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 622 nsew signal input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 623 nsew signal input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 624 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 625 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 626 nsew signal input
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 627 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 628 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 629 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 630 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 631 nsew signal tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 632 nsew signal tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 633 nsew signal tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 634 nsew signal tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 635 nsew signal tristate
rlabel metal4 s 576804 -1864 577404 705800 6 vccd1
port 636 nsew power bidirectional
rlabel metal4 s 540804 584916 541404 705800 6 vccd1.extra1
port 637 nsew power bidirectional
rlabel metal4 s 504804 584916 505404 705800 6 vccd1.extra2
port 638 nsew power bidirectional
rlabel metal4 s 468804 584916 469404 705800 6 vccd1.extra3
port 639 nsew power bidirectional
rlabel metal4 s 432804 584916 433404 705800 6 vccd1.extra4
port 640 nsew power bidirectional
rlabel metal4 s 396804 584916 397404 705800 6 vccd1.extra5
port 641 nsew power bidirectional
rlabel metal4 s 360804 584916 361404 705800 6 vccd1.extra6
port 642 nsew power bidirectional
rlabel metal4 s 324804 584916 325404 705800 6 vccd1.extra7
port 643 nsew power bidirectional
rlabel metal4 s 288804 356560 289404 705800 6 vccd1.extra8
port 644 nsew power bidirectional
rlabel metal4 s 252804 584916 253404 705800 6 vccd1.extra9
port 645 nsew power bidirectional
rlabel metal4 s 216804 584916 217404 705800 6 vccd1.extra10
port 646 nsew power bidirectional
rlabel metal4 s 180804 584916 181404 705800 6 vccd1.extra11
port 647 nsew power bidirectional
rlabel metal4 s 144804 584916 145404 705800 6 vccd1.extra12
port 648 nsew power bidirectional
rlabel metal4 s 108804 584916 109404 705800 6 vccd1.extra13
port 649 nsew power bidirectional
rlabel metal4 s 72804 584916 73404 705800 6 vccd1.extra14
port 650 nsew power bidirectional
rlabel metal4 s 36804 584916 37404 705800 6 vccd1.extra15
port 651 nsew power bidirectional
rlabel metal4 s 804 -1864 1404 705800 6 vccd1.extra16
port 652 nsew power bidirectional
rlabel metal4 s 585320 -924 585920 704860 6 vccd1.extra17
port 653 nsew power bidirectional
rlabel metal4 s -1996 -924 -1396 704860 4 vccd1.extra18
port 654 nsew power bidirectional
rlabel metal4 s 540804 274600 541404 382916 6 vccd1.extra19
port 655 nsew power bidirectional
rlabel metal4 s 504804 274600 505404 382916 6 vccd1.extra20
port 656 nsew power bidirectional
rlabel metal4 s 468804 274600 469404 382916 6 vccd1.extra21
port 657 nsew power bidirectional
rlabel metal4 s 432804 274600 433404 382916 6 vccd1.extra22
port 658 nsew power bidirectional
rlabel metal4 s 396804 274600 397404 382916 6 vccd1.extra23
port 659 nsew power bidirectional
rlabel metal4 s 360804 274600 361404 382916 6 vccd1.extra24
port 660 nsew power bidirectional
rlabel metal4 s 324804 274600 325404 382916 6 vccd1.extra25
port 661 nsew power bidirectional
rlabel metal4 s 252804 274600 253404 382916 6 vccd1.extra26
port 662 nsew power bidirectional
rlabel metal4 s 216804 274600 217404 382916 6 vccd1.extra27
port 663 nsew power bidirectional
rlabel metal4 s 180804 274600 181404 382916 6 vccd1.extra28
port 664 nsew power bidirectional
rlabel metal4 s 144804 274600 145404 382916 6 vccd1.extra29
port 665 nsew power bidirectional
rlabel metal4 s 108804 274600 109404 382916 6 vccd1.extra30
port 666 nsew power bidirectional
rlabel metal4 s 72804 274600 73404 382916 6 vccd1.extra31
port 667 nsew power bidirectional
rlabel metal4 s 36804 274600 37404 382916 6 vccd1.extra32
port 668 nsew power bidirectional
rlabel metal4 s 288804 -1864 289404 314560 6 vccd1.extra33
port 669 nsew power bidirectional
rlabel metal4 s 540804 -1864 541404 72600 6 vccd1.extra34
port 670 nsew power bidirectional
rlabel metal4 s 504804 -1864 505404 72600 6 vccd1.extra35
port 671 nsew power bidirectional
rlabel metal4 s 468804 -1864 469404 72600 6 vccd1.extra36
port 672 nsew power bidirectional
rlabel metal4 s 432804 -1864 433404 72600 6 vccd1.extra37
port 673 nsew power bidirectional
rlabel metal4 s 396804 -1864 397404 72600 6 vccd1.extra38
port 674 nsew power bidirectional
rlabel metal4 s 360804 -1864 361404 72600 6 vccd1.extra39
port 675 nsew power bidirectional
rlabel metal4 s 324804 -1864 325404 72600 6 vccd1.extra40
port 676 nsew power bidirectional
rlabel metal4 s 252804 -1864 253404 72600 6 vccd1.extra41
port 677 nsew power bidirectional
rlabel metal4 s 216804 -1864 217404 72600 6 vccd1.extra42
port 678 nsew power bidirectional
rlabel metal4 s 180804 -1864 181404 72600 6 vccd1.extra43
port 679 nsew power bidirectional
rlabel metal4 s 144804 -1864 145404 72600 6 vccd1.extra44
port 680 nsew power bidirectional
rlabel metal4 s 108804 -1864 109404 72600 6 vccd1.extra45
port 681 nsew power bidirectional
rlabel metal4 s 72804 -1864 73404 72600 6 vccd1.extra46
port 682 nsew power bidirectional
rlabel metal4 s 36804 -1864 37404 72600 6 vccd1.extra47
port 683 nsew power bidirectional
rlabel metal5 s -1996 704260 585920 704860 6 vccd1.extra48
port 684 nsew power bidirectional
rlabel metal5 s -2936 685876 586860 686476 6 vccd1.extra49
port 685 nsew power bidirectional
rlabel metal5 s -2936 649876 586860 650476 6 vccd1.extra50
port 686 nsew power bidirectional
rlabel metal5 s -2936 613876 586860 614476 6 vccd1.extra51
port 687 nsew power bidirectional
rlabel metal5 s -2936 577876 586860 578476 6 vccd1.extra52
port 688 nsew power bidirectional
rlabel metal5 s -2936 541876 586860 542476 6 vccd1.extra53
port 689 nsew power bidirectional
rlabel metal5 s -2936 505876 586860 506476 6 vccd1.extra54
port 690 nsew power bidirectional
rlabel metal5 s -2936 469876 586860 470476 6 vccd1.extra55
port 691 nsew power bidirectional
rlabel metal5 s -2936 433876 586860 434476 6 vccd1.extra56
port 692 nsew power bidirectional
rlabel metal5 s -2936 397876 586860 398476 6 vccd1.extra57
port 693 nsew power bidirectional
rlabel metal5 s -2936 361876 586860 362476 6 vccd1.extra58
port 694 nsew power bidirectional
rlabel metal5 s -2936 325876 586860 326476 6 vccd1.extra59
port 695 nsew power bidirectional
rlabel metal5 s -2936 289876 586860 290476 6 vccd1.extra60
port 696 nsew power bidirectional
rlabel metal5 s -2936 253876 586860 254476 6 vccd1.extra61
port 697 nsew power bidirectional
rlabel metal5 s -2936 217876 586860 218476 6 vccd1.extra62
port 698 nsew power bidirectional
rlabel metal5 s -2936 181876 586860 182476 6 vccd1.extra63
port 699 nsew power bidirectional
rlabel metal5 s -2936 145876 586860 146476 6 vccd1.extra64
port 700 nsew power bidirectional
rlabel metal5 s -2936 109876 586860 110476 6 vccd1.extra65
port 701 nsew power bidirectional
rlabel metal5 s -2936 73876 586860 74476 6 vccd1.extra66
port 702 nsew power bidirectional
rlabel metal5 s -2936 37876 586860 38476 6 vccd1.extra67
port 703 nsew power bidirectional
rlabel metal5 s -2936 1876 586860 2476 6 vccd1.extra68
port 704 nsew power bidirectional
rlabel metal5 s -1996 -924 585920 -324 8 vccd1.extra69
port 705 nsew power bidirectional
rlabel metal4 s 586260 -1864 586860 705800 6 vssd1
port 706 nsew ground bidirectional
rlabel metal4 s 558804 584916 559404 705800 6 vssd1.extra1
port 707 nsew ground bidirectional
rlabel metal4 s 522804 584916 523404 705800 6 vssd1.extra2
port 708 nsew ground bidirectional
rlabel metal4 s 486804 584916 487404 705800 6 vssd1.extra3
port 709 nsew ground bidirectional
rlabel metal4 s 450804 584916 451404 705800 6 vssd1.extra4
port 710 nsew ground bidirectional
rlabel metal4 s 414804 584916 415404 705800 6 vssd1.extra5
port 711 nsew ground bidirectional
rlabel metal4 s 378804 584916 379404 705800 6 vssd1.extra6
port 712 nsew ground bidirectional
rlabel metal4 s 342804 584916 343404 705800 6 vssd1.extra7
port 713 nsew ground bidirectional
rlabel metal4 s 306804 356560 307404 705800 6 vssd1.extra8
port 714 nsew ground bidirectional
rlabel metal4 s 270804 356560 271404 705800 6 vssd1.extra9
port 715 nsew ground bidirectional
rlabel metal4 s 234804 584916 235404 705800 6 vssd1.extra10
port 716 nsew ground bidirectional
rlabel metal4 s 198804 584916 199404 705800 6 vssd1.extra11
port 717 nsew ground bidirectional
rlabel metal4 s 162804 584916 163404 705800 6 vssd1.extra12
port 718 nsew ground bidirectional
rlabel metal4 s 126804 584916 127404 705800 6 vssd1.extra13
port 719 nsew ground bidirectional
rlabel metal4 s 90804 584916 91404 705800 6 vssd1.extra14
port 720 nsew ground bidirectional
rlabel metal4 s 54804 584916 55404 705800 6 vssd1.extra15
port 721 nsew ground bidirectional
rlabel metal4 s 18804 -1864 19404 705800 6 vssd1.extra16
port 722 nsew ground bidirectional
rlabel metal4 s -2936 -1864 -2336 705800 4 vssd1.extra17
port 723 nsew ground bidirectional
rlabel metal4 s 558804 274600 559404 382916 6 vssd1.extra18
port 724 nsew ground bidirectional
rlabel metal4 s 522804 274600 523404 382916 6 vssd1.extra19
port 725 nsew ground bidirectional
rlabel metal4 s 486804 274600 487404 382916 6 vssd1.extra20
port 726 nsew ground bidirectional
rlabel metal4 s 450804 274600 451404 382916 6 vssd1.extra21
port 727 nsew ground bidirectional
rlabel metal4 s 414804 274600 415404 382916 6 vssd1.extra22
port 728 nsew ground bidirectional
rlabel metal4 s 378804 274600 379404 382916 6 vssd1.extra23
port 729 nsew ground bidirectional
rlabel metal4 s 342804 274600 343404 382916 6 vssd1.extra24
port 730 nsew ground bidirectional
rlabel metal4 s 234804 274600 235404 382916 6 vssd1.extra25
port 731 nsew ground bidirectional
rlabel metal4 s 198804 274600 199404 382916 6 vssd1.extra26
port 732 nsew ground bidirectional
rlabel metal4 s 162804 274600 163404 382916 6 vssd1.extra27
port 733 nsew ground bidirectional
rlabel metal4 s 126804 274600 127404 382916 6 vssd1.extra28
port 734 nsew ground bidirectional
rlabel metal4 s 90804 274600 91404 382916 6 vssd1.extra29
port 735 nsew ground bidirectional
rlabel metal4 s 54804 274600 55404 382916 6 vssd1.extra30
port 736 nsew ground bidirectional
rlabel metal4 s 306804 -1864 307404 314560 6 vssd1.extra31
port 737 nsew ground bidirectional
rlabel metal4 s 270804 -1864 271404 314560 6 vssd1.extra32
port 738 nsew ground bidirectional
rlabel metal4 s 558804 -1864 559404 72600 6 vssd1.extra33
port 739 nsew ground bidirectional
rlabel metal4 s 522804 -1864 523404 72600 6 vssd1.extra34
port 740 nsew ground bidirectional
rlabel metal4 s 486804 -1864 487404 72600 6 vssd1.extra35
port 741 nsew ground bidirectional
rlabel metal4 s 450804 -1864 451404 72600 6 vssd1.extra36
port 742 nsew ground bidirectional
rlabel metal4 s 414804 -1864 415404 72600 6 vssd1.extra37
port 743 nsew ground bidirectional
rlabel metal4 s 378804 -1864 379404 72600 6 vssd1.extra38
port 744 nsew ground bidirectional
rlabel metal4 s 342804 -1864 343404 72600 6 vssd1.extra39
port 745 nsew ground bidirectional
rlabel metal4 s 234804 -1864 235404 72600 6 vssd1.extra40
port 746 nsew ground bidirectional
rlabel metal4 s 198804 -1864 199404 72600 6 vssd1.extra41
port 747 nsew ground bidirectional
rlabel metal4 s 162804 -1864 163404 72600 6 vssd1.extra42
port 748 nsew ground bidirectional
rlabel metal4 s 126804 -1864 127404 72600 6 vssd1.extra43
port 749 nsew ground bidirectional
rlabel metal4 s 90804 -1864 91404 72600 6 vssd1.extra44
port 750 nsew ground bidirectional
rlabel metal4 s 54804 -1864 55404 72600 6 vssd1.extra45
port 751 nsew ground bidirectional
rlabel metal5 s -2936 705200 586860 705800 6 vssd1.extra46
port 752 nsew ground bidirectional
rlabel metal5 s -2936 667876 586860 668476 6 vssd1.extra47
port 753 nsew ground bidirectional
rlabel metal5 s -2936 631876 586860 632476 6 vssd1.extra48
port 754 nsew ground bidirectional
rlabel metal5 s -2936 595876 586860 596476 6 vssd1.extra49
port 755 nsew ground bidirectional
rlabel metal5 s -2936 559876 586860 560476 6 vssd1.extra50
port 756 nsew ground bidirectional
rlabel metal5 s -2936 523876 586860 524476 6 vssd1.extra51
port 757 nsew ground bidirectional
rlabel metal5 s -2936 487876 586860 488476 6 vssd1.extra52
port 758 nsew ground bidirectional
rlabel metal5 s -2936 451876 586860 452476 6 vssd1.extra53
port 759 nsew ground bidirectional
rlabel metal5 s -2936 415876 586860 416476 6 vssd1.extra54
port 760 nsew ground bidirectional
rlabel metal5 s -2936 379876 586860 380476 6 vssd1.extra55
port 761 nsew ground bidirectional
rlabel metal5 s -2936 343876 586860 344476 6 vssd1.extra56
port 762 nsew ground bidirectional
rlabel metal5 s -2936 307876 586860 308476 6 vssd1.extra57
port 763 nsew ground bidirectional
rlabel metal5 s -2936 271876 586860 272476 6 vssd1.extra58
port 764 nsew ground bidirectional
rlabel metal5 s -2936 235876 586860 236476 6 vssd1.extra59
port 765 nsew ground bidirectional
rlabel metal5 s -2936 199876 586860 200476 6 vssd1.extra60
port 766 nsew ground bidirectional
rlabel metal5 s -2936 163876 586860 164476 6 vssd1.extra61
port 767 nsew ground bidirectional
rlabel metal5 s -2936 127876 586860 128476 6 vssd1.extra62
port 768 nsew ground bidirectional
rlabel metal5 s -2936 91876 586860 92476 6 vssd1.extra63
port 769 nsew ground bidirectional
rlabel metal5 s -2936 55876 586860 56476 6 vssd1.extra64
port 770 nsew ground bidirectional
rlabel metal5 s -2936 19876 586860 20476 6 vssd1.extra65
port 771 nsew ground bidirectional
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1.extra66
port 772 nsew ground bidirectional
rlabel metal4 s 587200 -2804 587800 706740 6 vccd2
port 773 nsew power bidirectional
rlabel metal4 s -3876 -2804 -3276 706740 4 vccd2.extra1
port 774 nsew power bidirectional
rlabel metal5 s -3876 706140 587800 706740 6 vccd2.extra2
port 775 nsew power bidirectional
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2.extra3
port 776 nsew power bidirectional
rlabel metal4 s 588140 -3744 588740 707680 6 vssd2
port 777 nsew ground bidirectional
rlabel metal4 s -4816 -3744 -4216 707680 4 vssd2.extra1
port 778 nsew ground bidirectional
rlabel metal5 s -4816 707080 588740 707680 6 vssd2.extra2
port 779 nsew ground bidirectional
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2.extra3
port 780 nsew ground bidirectional
rlabel metal4 s 589080 -4684 589680 708620 6 vdda1
port 781 nsew power bidirectional
rlabel metal4 s -5756 -4684 -5156 708620 4 vdda1.extra1
port 782 nsew power bidirectional
rlabel metal5 s -5756 708020 589680 708620 6 vdda1.extra2
port 783 nsew power bidirectional
rlabel metal5 s -5756 -4684 589680 -4084 8 vdda1.extra3
port 784 nsew power bidirectional
rlabel metal4 s 590020 -5624 590620 709560 6 vssa1
port 785 nsew ground bidirectional
rlabel metal4 s -6696 -5624 -6096 709560 4 vssa1.extra1
port 786 nsew ground bidirectional
rlabel metal5 s -6696 708960 590620 709560 6 vssa1.extra2
port 787 nsew ground bidirectional
rlabel metal5 s -6696 -5624 590620 -5024 8 vssa1.extra3
port 788 nsew ground bidirectional
rlabel metal4 s 590960 -6564 591560 710500 6 vdda2
port 789 nsew power bidirectional
rlabel metal4 s -7636 -6564 -7036 710500 4 vdda2.extra1
port 790 nsew power bidirectional
rlabel metal5 s -7636 709900 591560 710500 6 vdda2.extra2
port 791 nsew power bidirectional
rlabel metal5 s -7636 -6564 591560 -5964 8 vdda2.extra3
port 792 nsew power bidirectional
rlabel metal4 s 591900 -7504 592500 711440 6 vssa2
port 793 nsew ground bidirectional
rlabel metal4 s -8576 -7504 -7976 711440 4 vssa2.extra1
port 794 nsew ground bidirectional
rlabel metal5 s -8576 710840 592500 711440 6 vssa2.extra2
port 795 nsew ground bidirectional
rlabel metal5 s -8576 -7504 592500 -6904 8 vssa2.extra3
port 796 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>

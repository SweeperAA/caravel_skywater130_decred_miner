magic
tech sky130A
magscale 1 2
timestamp 1608091038
<< locali >>
rect 340061 586483 340095 586585
rect 233985 586143 234019 586313
rect 319453 586211 319487 586449
rect 329665 586211 329699 586449
rect 348893 586483 348927 586585
rect 381277 586483 381311 586585
rect 329757 586279 329791 586449
rect 369501 586279 369535 586381
rect 379713 586279 379747 586449
rect 391489 586415 391523 586585
rect 401885 586483 401919 586585
rect 412097 586415 412131 586585
rect 422493 586483 422527 586585
rect 432705 586415 432739 586585
rect 443101 586483 443135 586585
rect 453313 586415 453347 586585
rect 463709 586483 463743 586585
rect 473921 586415 473955 586585
rect 394467 586381 394525 586415
rect 415075 586381 415133 586415
rect 435683 586381 435741 586415
rect 456291 586381 456349 586415
rect 476899 586381 476957 586415
rect 198749 585939 198783 586109
rect 244381 585939 244415 586109
rect 254593 585939 254627 586109
rect 314301 494615 314335 504849
rect 314301 474011 314335 484245
rect 314301 453407 314335 463641
rect 314393 425391 314427 432701
rect 269865 340051 269899 350285
rect 272901 340051 272935 343009
rect 270049 297415 270083 309077
rect 269865 287079 269899 293301
rect 188445 276403 188479 276505
rect 177313 276131 177347 276233
rect 195805 276199 195839 276301
rect 204637 276063 204671 276301
rect 214941 276267 214975 276437
rect 225153 276267 225187 276437
rect 257629 276199 257663 276437
rect 267841 276199 267875 276437
rect 278145 276403 278179 276641
rect 288541 276199 288575 276573
rect 368029 276199 368063 276369
rect 209697 276063 209731 276165
rect 306205 275927 306239 276165
rect 316417 275927 316451 276165
rect 326813 275927 326847 276165
rect 337025 275927 337059 276165
rect 347421 275995 347455 276165
rect 378241 276199 378275 276369
rect 388637 276199 388671 276369
rect 394525 276267 394559 276369
rect 404829 276199 404863 276437
rect 453405 276335 453439 276437
rect 435683 276301 435741 276335
rect 357633 275995 357667 276165
rect 270141 144279 270175 152881
rect 270141 120751 270175 130985
rect 269807 72097 270049 72131
<< viali >>
rect 340061 586585 340095 586619
rect 319453 586449 319487 586483
rect 233985 586313 234019 586347
rect 319453 586177 319487 586211
rect 329665 586449 329699 586483
rect 329757 586449 329791 586483
rect 340061 586449 340095 586483
rect 348893 586585 348927 586619
rect 381277 586585 381311 586619
rect 348893 586449 348927 586483
rect 379713 586449 379747 586483
rect 381277 586449 381311 586483
rect 391489 586585 391523 586619
rect 329757 586245 329791 586279
rect 369501 586381 369535 586415
rect 369501 586245 369535 586279
rect 401885 586585 401919 586619
rect 401885 586449 401919 586483
rect 412097 586585 412131 586619
rect 422493 586585 422527 586619
rect 422493 586449 422527 586483
rect 432705 586585 432739 586619
rect 443101 586585 443135 586619
rect 443101 586449 443135 586483
rect 453313 586585 453347 586619
rect 463709 586585 463743 586619
rect 463709 586449 463743 586483
rect 473921 586585 473955 586619
rect 391489 586381 391523 586415
rect 394433 586381 394467 586415
rect 394525 586381 394559 586415
rect 412097 586381 412131 586415
rect 415041 586381 415075 586415
rect 415133 586381 415167 586415
rect 432705 586381 432739 586415
rect 435649 586381 435683 586415
rect 435741 586381 435775 586415
rect 453313 586381 453347 586415
rect 456257 586381 456291 586415
rect 456349 586381 456383 586415
rect 473921 586381 473955 586415
rect 476865 586381 476899 586415
rect 476957 586381 476991 586415
rect 379713 586245 379747 586279
rect 329665 586177 329699 586211
rect 198749 586109 198783 586143
rect 233985 586109 234019 586143
rect 244381 586109 244415 586143
rect 198749 585905 198783 585939
rect 244381 585905 244415 585939
rect 254593 586109 254627 586143
rect 254593 585905 254627 585939
rect 314301 504849 314335 504883
rect 314301 494581 314335 494615
rect 314301 484245 314335 484279
rect 314301 473977 314335 474011
rect 314301 463641 314335 463675
rect 314301 453373 314335 453407
rect 314393 432701 314427 432735
rect 314393 425357 314427 425391
rect 269865 350285 269899 350319
rect 269865 340017 269899 340051
rect 272901 343009 272935 343043
rect 272901 340017 272935 340051
rect 270049 309077 270083 309111
rect 270049 297381 270083 297415
rect 269865 293301 269899 293335
rect 269865 287045 269899 287079
rect 278145 276641 278179 276675
rect 188445 276505 188479 276539
rect 188445 276369 188479 276403
rect 214941 276437 214975 276471
rect 195805 276301 195839 276335
rect 177313 276233 177347 276267
rect 195805 276165 195839 276199
rect 204637 276301 204671 276335
rect 177313 276097 177347 276131
rect 214941 276233 214975 276267
rect 225153 276437 225187 276471
rect 225153 276233 225187 276267
rect 257629 276437 257663 276471
rect 204637 276029 204671 276063
rect 209697 276165 209731 276199
rect 257629 276165 257663 276199
rect 267841 276437 267875 276471
rect 278145 276369 278179 276403
rect 288541 276573 288575 276607
rect 267841 276165 267875 276199
rect 404829 276437 404863 276471
rect 368029 276369 368063 276403
rect 288541 276165 288575 276199
rect 306205 276165 306239 276199
rect 209697 276029 209731 276063
rect 306205 275893 306239 275927
rect 316417 276165 316451 276199
rect 316417 275893 316451 275927
rect 326813 276165 326847 276199
rect 326813 275893 326847 275927
rect 337025 276165 337059 276199
rect 347421 276165 347455 276199
rect 347421 275961 347455 275995
rect 357633 276165 357667 276199
rect 368029 276165 368063 276199
rect 378241 276369 378275 276403
rect 378241 276165 378275 276199
rect 388637 276369 388671 276403
rect 394525 276369 394559 276403
rect 394525 276233 394559 276267
rect 388637 276165 388671 276199
rect 453405 276437 453439 276471
rect 435649 276301 435683 276335
rect 435741 276301 435775 276335
rect 453405 276301 453439 276335
rect 404829 276165 404863 276199
rect 357633 275961 357667 275995
rect 337025 275893 337059 275927
rect 270141 152881 270175 152915
rect 270141 144245 270175 144279
rect 270141 130985 270175 131019
rect 270141 120717 270175 120751
rect 269773 72097 269807 72131
rect 270049 72097 270083 72131
<< metal1 >>
rect 8018 700612 8024 700664
rect 8076 700652 8082 700664
rect 8202 700652 8208 700664
rect 8076 700624 8208 700652
rect 8076 700612 8082 700624
rect 8202 700612 8208 700624
rect 8260 700652 8266 700664
rect 72970 700652 72976 700664
rect 8260 700624 72976 700652
rect 8260 700612 8266 700624
rect 72970 700612 72976 700624
rect 73028 700652 73034 700664
rect 137830 700652 137836 700664
rect 73028 700624 137836 700652
rect 73028 700612 73034 700624
rect 137830 700612 137836 700624
rect 137888 700652 137894 700664
rect 202782 700652 202788 700664
rect 137888 700624 202788 700652
rect 137888 700612 137894 700624
rect 202782 700612 202788 700624
rect 202840 700652 202846 700664
rect 267642 700652 267648 700664
rect 202840 700624 267648 700652
rect 202840 700612 202846 700624
rect 267642 700612 267648 700624
rect 267700 700652 267706 700664
rect 273806 700652 273812 700664
rect 267700 700624 273812 700652
rect 267700 700612 267706 700624
rect 273806 700612 273812 700624
rect 273864 700612 273870 700664
rect 332502 700612 332508 700664
rect 332560 700652 332566 700664
rect 397454 700652 397460 700664
rect 332560 700624 397460 700652
rect 332560 700612 332566 700624
rect 397454 700612 397460 700624
rect 397512 700652 397518 700664
rect 462314 700652 462320 700664
rect 397512 700624 462320 700652
rect 397512 700612 397518 700624
rect 462314 700612 462320 700624
rect 462372 700652 462378 700664
rect 527174 700652 527180 700664
rect 462372 700624 527180 700652
rect 462372 700612 462378 700624
rect 527174 700612 527180 700624
rect 527232 700612 527238 700664
rect 272978 700068 272984 700120
rect 273036 700108 273042 700120
rect 283834 700108 283840 700120
rect 273036 700080 283840 700108
rect 273036 700068 273042 700080
rect 283834 700068 283840 700080
rect 283892 700068 283898 700120
rect 273070 700000 273076 700052
rect 273128 700040 273134 700052
rect 364978 700040 364984 700052
rect 273128 700012 364984 700040
rect 273128 700000 273134 700012
rect 364978 700000 364984 700012
rect 365036 700000 365042 700052
rect 270678 699932 270684 699984
rect 270736 699972 270742 699984
rect 429838 699972 429844 699984
rect 270736 699944 429844 699972
rect 270736 699932 270742 699944
rect 429838 699932 429844 699944
rect 429896 699932 429902 699984
rect 527174 699932 527180 699984
rect 527232 699972 527238 699984
rect 579890 699972 579896 699984
rect 527232 699944 579896 699972
rect 527232 699932 527238 699944
rect 579890 699932 579896 699944
rect 579948 699932 579954 699984
rect 154114 699864 154120 699916
rect 154172 699904 154178 699916
rect 268562 699904 268568 699916
rect 154172 699876 268568 699904
rect 154172 699864 154178 699876
rect 268562 699864 268568 699876
rect 268620 699864 268626 699916
rect 270770 699864 270776 699916
rect 270828 699904 270834 699916
rect 559650 699904 559656 699916
rect 270828 699876 559656 699904
rect 270828 699864 270834 699876
rect 559650 699864 559656 699876
rect 559708 699864 559714 699916
rect 2958 653488 2964 653540
rect 3016 653528 3022 653540
rect 8018 653528 8024 653540
rect 3016 653500 8024 653528
rect 3016 653488 3022 653500
rect 8018 653488 8024 653500
rect 8076 653488 8082 653540
rect 270494 627104 270500 627156
rect 270552 627144 270558 627156
rect 578786 627144 578792 627156
rect 270552 627116 578792 627144
rect 270552 627104 270558 627116
rect 578786 627104 578792 627116
rect 578844 627104 578850 627156
rect 340049 586619 340107 586625
rect 340049 586585 340061 586619
rect 340095 586616 340107 586619
rect 348881 586619 348939 586625
rect 348881 586616 348893 586619
rect 340095 586588 348893 586616
rect 340095 586585 340107 586588
rect 340049 586579 340107 586585
rect 348881 586585 348893 586588
rect 348927 586585 348939 586619
rect 348881 586579 348939 586585
rect 381265 586619 381323 586625
rect 381265 586585 381277 586619
rect 381311 586616 381323 586619
rect 391477 586619 391535 586625
rect 391477 586616 391489 586619
rect 381311 586588 391489 586616
rect 381311 586585 381323 586588
rect 381265 586579 381323 586585
rect 391477 586585 391489 586588
rect 391523 586585 391535 586619
rect 391477 586579 391535 586585
rect 401873 586619 401931 586625
rect 401873 586585 401885 586619
rect 401919 586616 401931 586619
rect 412085 586619 412143 586625
rect 412085 586616 412097 586619
rect 401919 586588 412097 586616
rect 401919 586585 401931 586588
rect 401873 586579 401931 586585
rect 412085 586585 412097 586588
rect 412131 586585 412143 586619
rect 412085 586579 412143 586585
rect 422481 586619 422539 586625
rect 422481 586585 422493 586619
rect 422527 586616 422539 586619
rect 432693 586619 432751 586625
rect 432693 586616 432705 586619
rect 422527 586588 432705 586616
rect 422527 586585 422539 586588
rect 422481 586579 422539 586585
rect 432693 586585 432705 586588
rect 432739 586585 432751 586619
rect 432693 586579 432751 586585
rect 443089 586619 443147 586625
rect 443089 586585 443101 586619
rect 443135 586616 443147 586619
rect 453301 586619 453359 586625
rect 453301 586616 453313 586619
rect 443135 586588 453313 586616
rect 443135 586585 443147 586588
rect 443089 586579 443147 586585
rect 453301 586585 453313 586588
rect 453347 586585 453359 586619
rect 453301 586579 453359 586585
rect 463697 586619 463755 586625
rect 463697 586585 463709 586619
rect 463743 586616 463755 586619
rect 473909 586619 473967 586625
rect 473909 586616 473921 586619
rect 463743 586588 473921 586616
rect 463743 586585 463755 586588
rect 463697 586579 463755 586585
rect 473909 586585 473921 586588
rect 473955 586585 473967 586619
rect 473909 586579 473967 586585
rect 49602 586440 49608 586492
rect 49660 586480 49666 586492
rect 307570 586480 307576 586492
rect 49660 586452 307576 586480
rect 49660 586440 49666 586452
rect 307570 586440 307576 586452
rect 307628 586440 307634 586492
rect 319441 586483 319499 586489
rect 319441 586449 319453 586483
rect 319487 586480 319499 586483
rect 329653 586483 329711 586489
rect 329653 586480 329665 586483
rect 319487 586452 329665 586480
rect 319487 586449 319499 586452
rect 319441 586443 319499 586449
rect 329653 586449 329665 586452
rect 329699 586449 329711 586483
rect 329653 586443 329711 586449
rect 329745 586483 329803 586489
rect 329745 586449 329757 586483
rect 329791 586480 329803 586483
rect 340049 586483 340107 586489
rect 340049 586480 340061 586483
rect 329791 586452 340061 586480
rect 329791 586449 329803 586452
rect 329745 586443 329803 586449
rect 340049 586449 340061 586452
rect 340095 586449 340107 586483
rect 340049 586443 340107 586449
rect 348881 586483 348939 586489
rect 348881 586449 348893 586483
rect 348927 586480 348939 586483
rect 379701 586483 379759 586489
rect 348927 586452 359136 586480
rect 348927 586449 348939 586452
rect 348881 586443 348939 586449
rect 73522 586372 73528 586424
rect 73580 586412 73586 586424
rect 289446 586412 289452 586424
rect 73580 586384 289452 586412
rect 73580 586372 73586 586384
rect 289446 586372 289452 586384
rect 289504 586372 289510 586424
rect 359108 586412 359136 586452
rect 379701 586449 379713 586483
rect 379747 586480 379759 586483
rect 381265 586483 381323 586489
rect 381265 586480 381277 586483
rect 379747 586452 381277 586480
rect 379747 586449 379759 586452
rect 379701 586443 379759 586449
rect 381265 586449 381277 586452
rect 381311 586449 381323 586483
rect 401873 586483 401931 586489
rect 401873 586480 401885 586483
rect 381265 586443 381323 586449
rect 396644 586452 401885 586480
rect 369489 586415 369547 586421
rect 369489 586412 369501 586415
rect 359108 586384 369501 586412
rect 369489 586381 369501 586384
rect 369535 586381 369547 586415
rect 369489 586375 369547 586381
rect 391477 586415 391535 586421
rect 391477 586381 391489 586415
rect 391523 586412 391535 586415
rect 394421 586415 394479 586421
rect 394421 586412 394433 586415
rect 391523 586384 394433 586412
rect 391523 586381 391535 586384
rect 391477 586375 391535 586381
rect 394421 586381 394433 586384
rect 394467 586381 394479 586415
rect 394421 586375 394479 586381
rect 394513 586415 394571 586421
rect 394513 586381 394525 586415
rect 394559 586412 394571 586415
rect 396644 586412 396672 586452
rect 401873 586449 401885 586452
rect 401919 586449 401931 586483
rect 422481 586483 422539 586489
rect 422481 586480 422493 586483
rect 401873 586443 401931 586449
rect 417252 586452 422493 586480
rect 394559 586384 396672 586412
rect 412085 586415 412143 586421
rect 394559 586381 394571 586384
rect 394513 586375 394571 586381
rect 412085 586381 412097 586415
rect 412131 586412 412143 586415
rect 415029 586415 415087 586421
rect 415029 586412 415041 586415
rect 412131 586384 415041 586412
rect 412131 586381 412143 586384
rect 412085 586375 412143 586381
rect 415029 586381 415041 586384
rect 415075 586381 415087 586415
rect 415029 586375 415087 586381
rect 415121 586415 415179 586421
rect 415121 586381 415133 586415
rect 415167 586412 415179 586415
rect 417252 586412 417280 586452
rect 422481 586449 422493 586452
rect 422527 586449 422539 586483
rect 443089 586483 443147 586489
rect 443089 586480 443101 586483
rect 422481 586443 422539 586449
rect 437860 586452 443101 586480
rect 415167 586384 417280 586412
rect 432693 586415 432751 586421
rect 415167 586381 415179 586384
rect 415121 586375 415179 586381
rect 432693 586381 432705 586415
rect 432739 586412 432751 586415
rect 435637 586415 435695 586421
rect 435637 586412 435649 586415
rect 432739 586384 435649 586412
rect 432739 586381 432751 586384
rect 432693 586375 432751 586381
rect 435637 586381 435649 586384
rect 435683 586381 435695 586415
rect 435637 586375 435695 586381
rect 435729 586415 435787 586421
rect 435729 586381 435741 586415
rect 435775 586412 435787 586415
rect 437860 586412 437888 586452
rect 443089 586449 443101 586452
rect 443135 586449 443147 586483
rect 463697 586483 463755 586489
rect 463697 586480 463709 586483
rect 443089 586443 443147 586449
rect 458468 586452 463709 586480
rect 435775 586384 437888 586412
rect 453301 586415 453359 586421
rect 435775 586381 435787 586384
rect 435729 586375 435787 586381
rect 453301 586381 453313 586415
rect 453347 586412 453359 586415
rect 456245 586415 456303 586421
rect 456245 586412 456257 586415
rect 453347 586384 456257 586412
rect 453347 586381 453359 586384
rect 453301 586375 453359 586381
rect 456245 586381 456257 586384
rect 456291 586381 456303 586415
rect 456245 586375 456303 586381
rect 456337 586415 456395 586421
rect 456337 586381 456349 586415
rect 456383 586412 456395 586415
rect 458468 586412 458496 586452
rect 463697 586449 463709 586452
rect 463743 586449 463755 586483
rect 485774 586480 485780 586492
rect 463697 586443 463755 586449
rect 479076 586452 485780 586480
rect 456383 586384 458496 586412
rect 473909 586415 473967 586421
rect 456383 586381 456395 586384
rect 456337 586375 456395 586381
rect 473909 586381 473921 586415
rect 473955 586412 473967 586415
rect 476853 586415 476911 586421
rect 476853 586412 476865 586415
rect 473955 586384 476865 586412
rect 473955 586381 473967 586384
rect 473909 586375 473967 586381
rect 476853 586381 476865 586384
rect 476899 586381 476911 586415
rect 476853 586375 476911 586381
rect 476945 586415 477003 586421
rect 476945 586381 476957 586415
rect 476991 586412 477003 586415
rect 479076 586412 479104 586452
rect 485774 586440 485780 586452
rect 485832 586440 485838 586492
rect 476991 586384 479104 586412
rect 476991 586381 477003 586384
rect 476945 586375 477003 586381
rect 219342 586304 219348 586356
rect 219400 586344 219406 586356
rect 233973 586347 234031 586353
rect 233973 586344 233985 586347
rect 219400 586316 233985 586344
rect 219400 586304 219406 586316
rect 233973 586313 233985 586316
rect 234019 586313 234031 586347
rect 233973 586307 234031 586313
rect 242066 586304 242072 586356
rect 242124 586344 242130 586356
rect 293586 586344 293592 586356
rect 242124 586316 293592 586344
rect 242124 586304 242130 586316
rect 293586 586304 293592 586316
rect 293644 586304 293650 586356
rect 169754 586236 169760 586288
rect 169812 586276 169818 586288
rect 298646 586276 298652 586288
rect 169812 586248 298652 586276
rect 169812 586236 169818 586248
rect 298646 586236 298652 586248
rect 298704 586236 298710 586288
rect 329745 586279 329803 586285
rect 329745 586276 329757 586279
rect 329668 586248 329757 586276
rect 329668 586217 329696 586248
rect 329745 586245 329757 586248
rect 329791 586245 329803 586279
rect 329745 586239 329803 586245
rect 369489 586279 369547 586285
rect 369489 586245 369501 586279
rect 369535 586276 369547 586279
rect 379701 586279 379759 586285
rect 379701 586276 379713 586279
rect 369535 586248 379713 586276
rect 369535 586245 369547 586248
rect 369489 586239 369547 586245
rect 379701 586245 379713 586248
rect 379747 586245 379759 586279
rect 379701 586239 379759 586245
rect 319441 586211 319499 586217
rect 319441 586208 319453 586211
rect 270420 586180 319453 586208
rect 270420 586152 270448 586180
rect 319441 586177 319453 586180
rect 319487 586177 319499 586211
rect 319441 586171 319499 586177
rect 329653 586211 329711 586217
rect 329653 586177 329665 586211
rect 329699 586177 329711 586211
rect 329653 586171 329711 586177
rect 193858 586100 193864 586152
rect 193916 586140 193922 586152
rect 198737 586143 198795 586149
rect 198737 586140 198749 586143
rect 193916 586112 198749 586140
rect 193916 586100 193922 586112
rect 198737 586109 198749 586112
rect 198783 586109 198795 586143
rect 198737 586103 198795 586109
rect 233973 586143 234031 586149
rect 233973 586109 233985 586143
rect 234019 586140 234031 586143
rect 244369 586143 244427 586149
rect 244369 586140 244381 586143
rect 234019 586112 244381 586140
rect 234019 586109 234031 586112
rect 233973 586103 234031 586109
rect 244369 586109 244381 586112
rect 244415 586109 244427 586143
rect 244369 586103 244427 586109
rect 254581 586143 254639 586149
rect 254581 586109 254593 586143
rect 254627 586140 254639 586143
rect 270402 586140 270408 586152
rect 254627 586112 270408 586140
rect 254627 586109 254639 586112
rect 254581 586103 254639 586109
rect 270402 586100 270408 586112
rect 270460 586100 270466 586152
rect 270586 586100 270592 586152
rect 270644 586140 270650 586152
rect 509878 586140 509884 586152
rect 270644 586112 509884 586140
rect 270644 586100 270650 586112
rect 509878 586100 509884 586112
rect 509936 586100 509942 586152
rect 145834 586032 145840 586084
rect 145892 586072 145898 586084
rect 284754 586072 284760 586084
rect 145892 586044 284760 586072
rect 145892 586032 145898 586044
rect 284754 586032 284760 586044
rect 284812 586032 284818 586084
rect 293586 586032 293592 586084
rect 293644 586072 293650 586084
rect 533982 586072 533988 586084
rect 293644 586044 533988 586072
rect 293644 586032 293650 586044
rect 533982 586032 533988 586044
rect 534040 586032 534046 586084
rect 217962 585964 217968 586016
rect 218020 586004 218026 586016
rect 270586 586004 270592 586016
rect 218020 585976 270592 586004
rect 218020 585964 218026 585976
rect 270586 585964 270592 585976
rect 270644 585964 270650 586016
rect 300210 585964 300216 586016
rect 300268 586004 300274 586016
rect 437750 586004 437756 586016
rect 300268 585976 437756 586004
rect 300268 585964 300274 585976
rect 437750 585964 437756 585976
rect 437808 585964 437814 586016
rect 198737 585939 198795 585945
rect 198737 585905 198749 585939
rect 198783 585936 198795 585939
rect 219342 585936 219348 585948
rect 198783 585908 219348 585936
rect 198783 585905 198795 585908
rect 198737 585899 198795 585905
rect 219342 585896 219348 585908
rect 219400 585896 219406 585948
rect 244369 585939 244427 585945
rect 244369 585905 244381 585939
rect 244415 585936 244427 585939
rect 254581 585939 254639 585945
rect 254581 585936 254593 585939
rect 244415 585908 254593 585936
rect 244415 585905 244427 585908
rect 244369 585899 244427 585905
rect 254581 585905 254593 585908
rect 254627 585905 254639 585939
rect 254581 585899 254639 585905
rect 265986 585896 265992 585948
rect 266044 585936 266050 585948
rect 289170 585936 289176 585948
rect 266044 585908 289176 585936
rect 266044 585896 266050 585908
rect 289170 585896 289176 585908
rect 289228 585936 289234 585948
rect 557902 585936 557908 585948
rect 289228 585908 557908 585936
rect 289228 585896 289234 585908
rect 557902 585896 557908 585908
rect 557960 585896 557966 585948
rect 24854 582428 24860 582480
rect 24912 582468 24918 582480
rect 314378 582468 314384 582480
rect 24912 582440 314384 582468
rect 24912 582428 24918 582440
rect 314378 582428 314384 582440
rect 314436 582428 314442 582480
rect 26510 582360 26516 582412
rect 26568 582400 26574 582412
rect 267090 582400 267096 582412
rect 26568 582372 267096 582400
rect 26568 582360 26574 582372
rect 267090 582360 267096 582372
rect 267148 582360 267154 582412
rect 27246 582292 27252 582344
rect 27304 582332 27310 582344
rect 276658 582332 276664 582344
rect 27304 582304 276664 582332
rect 27304 582292 27310 582304
rect 276658 582292 276664 582304
rect 276716 582292 276722 582344
rect 319438 582292 319444 582344
rect 319496 582332 319502 582344
rect 558730 582332 558736 582344
rect 319496 582304 558736 582332
rect 319496 582292 319502 582304
rect 558730 582292 558736 582304
rect 558788 582292 558794 582344
rect 313458 582224 313464 582276
rect 313516 582264 313522 582276
rect 560846 582264 560852 582276
rect 313516 582236 560852 582264
rect 313516 582224 313522 582236
rect 560846 582224 560852 582236
rect 560904 582224 560910 582276
rect 276658 580660 276664 580712
rect 276716 580700 276722 580712
rect 315390 580700 315396 580712
rect 276716 580672 315396 580700
rect 276716 580660 276722 580672
rect 315390 580660 315396 580672
rect 315448 580660 315454 580712
rect 558546 579980 558552 580032
rect 558604 580020 558610 580032
rect 578786 580020 578792 580032
rect 558604 579992 578792 580020
rect 558604 579980 558610 579992
rect 578786 579980 578792 579992
rect 578844 579980 578850 580032
rect 317966 578484 317972 578536
rect 318024 578524 318030 578536
rect 319438 578524 319444 578536
rect 318024 578496 319444 578524
rect 318024 578484 318030 578496
rect 319438 578484 319444 578496
rect 319496 578484 319502 578536
rect 267090 575492 267096 575544
rect 267148 575532 267154 575544
rect 271874 575532 271880 575544
rect 267148 575504 271880 575532
rect 267148 575492 267154 575504
rect 271874 575492 271880 575504
rect 271932 575492 271938 575544
rect 26510 574104 26516 574116
rect 25056 574076 26516 574104
rect 24946 573996 24952 574048
rect 25004 574036 25010 574048
rect 25056 574036 25084 574076
rect 26510 574064 26516 574076
rect 26568 574064 26574 574116
rect 317966 574104 317972 574116
rect 310624 574076 317972 574104
rect 25004 574008 25084 574036
rect 25004 573996 25010 574008
rect 309134 573996 309140 574048
rect 309192 574036 309198 574048
rect 310624 574036 310652 574076
rect 317966 574064 317972 574076
rect 318024 574064 318030 574116
rect 309192 574008 310652 574036
rect 309192 573996 309198 574008
rect 305362 571820 305368 571872
rect 305420 571860 305426 571872
rect 309134 571860 309140 571872
rect 305420 571832 309140 571860
rect 305420 571820 305426 571832
rect 309134 571820 309140 571832
rect 309192 571820 309198 571872
rect 271874 571208 271880 571260
rect 271932 571248 271938 571260
rect 271932 571220 273852 571248
rect 271932 571208 271938 571220
rect 273824 571112 273852 571220
rect 276566 571112 276572 571124
rect 273824 571084 276572 571112
rect 276566 571072 276572 571084
rect 276624 571072 276630 571124
rect 276566 566652 276572 566704
rect 276624 566692 276630 566704
rect 279234 566692 279240 566704
rect 276624 566664 279240 566692
rect 276624 566652 276630 566664
rect 279234 566652 279240 566664
rect 279292 566652 279298 566704
rect 314102 565224 314108 565276
rect 314160 565264 314166 565276
rect 314378 565264 314384 565276
rect 314160 565236 314384 565264
rect 314160 565224 314166 565236
rect 314378 565224 314384 565236
rect 314436 565224 314442 565276
rect 279234 560056 279240 560108
rect 279292 560096 279298 560108
rect 280338 560096 280344 560108
rect 279292 560068 280344 560096
rect 279292 560056 279298 560068
rect 280338 560056 280344 560068
rect 280396 560056 280402 560108
rect 305362 557920 305368 557932
rect 303264 557892 305368 557920
rect 301682 557812 301688 557864
rect 301740 557852 301746 557864
rect 303264 557852 303292 557892
rect 305362 557880 305368 557892
rect 305420 557880 305426 557932
rect 301740 557824 303292 557852
rect 301740 557812 301746 557824
rect 299566 554344 299572 554396
rect 299624 554384 299630 554396
rect 301682 554384 301688 554396
rect 299624 554356 301688 554384
rect 299624 554344 299630 554356
rect 301682 554344 301688 554356
rect 301740 554344 301746 554396
rect 297358 552032 297364 552084
rect 297416 552072 297422 552084
rect 299566 552072 299572 552084
rect 297416 552044 299572 552072
rect 297416 552032 297422 552044
rect 299566 552032 299572 552044
rect 299624 552032 299630 552084
rect 268286 548972 268292 549024
rect 268344 549012 268350 549024
rect 313458 549012 313464 549024
rect 268344 548984 313464 549012
rect 268344 548972 268350 548984
rect 313458 548972 313464 548984
rect 313516 548972 313522 549024
rect 313458 547612 313464 547664
rect 313516 547652 313522 547664
rect 313918 547652 313924 547664
rect 313516 547624 313924 547652
rect 313516 547612 313522 547624
rect 313918 547612 313924 547624
rect 313976 547612 313982 547664
rect 314194 544824 314200 544876
rect 314252 544864 314258 544876
rect 315850 544864 315856 544876
rect 314252 544836 315856 544864
rect 314252 544824 314258 544836
rect 315850 544824 315856 544836
rect 315908 544824 315914 544876
rect 295886 543736 295892 543788
rect 295944 543776 295950 543788
rect 297358 543776 297364 543788
rect 295944 543748 297364 543776
rect 295944 543736 295950 543748
rect 297358 543736 297364 543748
rect 297416 543736 297422 543788
rect 280338 538704 280344 538756
rect 280396 538744 280402 538756
rect 282178 538744 282184 538756
rect 280396 538716 282184 538744
rect 280396 538704 280402 538716
rect 282178 538704 282184 538716
rect 282236 538704 282242 538756
rect 294414 538024 294420 538076
rect 294472 538064 294478 538076
rect 295886 538064 295892 538076
rect 294472 538036 295892 538064
rect 294472 538024 294478 538036
rect 295886 538024 295892 538036
rect 295944 538024 295950 538076
rect 282178 535032 282184 535084
rect 282236 535072 282242 535084
rect 288526 535072 288532 535084
rect 282236 535044 288532 535072
rect 282236 535032 282242 535044
rect 288526 535032 288532 535044
rect 288584 535032 288590 535084
rect 288526 533944 288532 533996
rect 288584 533984 288590 533996
rect 289998 533984 290004 533996
rect 288584 533956 290004 533984
rect 288584 533944 288590 533956
rect 289998 533944 290004 533956
rect 290056 533944 290062 533996
rect 291378 533672 291384 533724
rect 291436 533712 291442 533724
rect 294414 533712 294420 533724
rect 291436 533684 294420 533712
rect 291436 533672 291442 533684
rect 294414 533672 294420 533684
rect 294472 533672 294478 533724
rect 558638 532856 558644 532908
rect 558696 532896 558702 532908
rect 578786 532896 578792 532908
rect 558696 532868 578792 532896
rect 558696 532856 558702 532868
rect 578786 532856 578792 532868
rect 578844 532856 578850 532908
rect 289262 528436 289268 528488
rect 289320 528476 289326 528488
rect 291378 528476 291384 528488
rect 289320 528448 291384 528476
rect 289320 528436 289326 528448
rect 291378 528436 291384 528448
rect 291436 528436 291442 528488
rect 289998 526940 290004 526992
rect 290056 526980 290062 526992
rect 292758 526980 292764 526992
rect 290056 526952 292764 526980
rect 290056 526940 290062 526952
rect 292758 526940 292764 526952
rect 292816 526940 292822 526992
rect 292758 524016 292764 524068
rect 292816 524056 292822 524068
rect 292816 524028 292988 524056
rect 292816 524016 292822 524028
rect 292960 523988 292988 524028
rect 295518 523988 295524 524000
rect 292960 523960 295524 523988
rect 295518 523948 295524 523960
rect 295576 523948 295582 524000
rect 287054 523200 287060 523252
rect 287112 523240 287118 523252
rect 289262 523240 289268 523252
rect 287112 523212 289268 523240
rect 287112 523200 287118 523212
rect 289262 523200 289268 523212
rect 289320 523200 289326 523252
rect 295518 521024 295524 521076
rect 295576 521064 295582 521076
rect 298462 521064 298468 521076
rect 295576 521036 298468 521064
rect 295576 521024 295582 521036
rect 298462 521024 298468 521036
rect 298520 521024 298526 521076
rect 284110 516672 284116 516724
rect 284168 516712 284174 516724
rect 286962 516712 286968 516724
rect 284168 516684 286968 516712
rect 284168 516672 284174 516684
rect 286962 516672 286968 516684
rect 287020 516672 287026 516724
rect 298462 516672 298468 516724
rect 298520 516712 298526 516724
rect 301774 516712 301780 516724
rect 298520 516684 301780 516712
rect 298520 516672 298526 516684
rect 301774 516672 301780 516684
rect 301832 516672 301838 516724
rect 283282 515176 283288 515228
rect 283340 515216 283346 515228
rect 284110 515216 284116 515228
rect 283340 515188 284116 515216
rect 283340 515176 283346 515188
rect 284110 515176 284116 515188
rect 284168 515176 284174 515228
rect 558730 515108 558736 515160
rect 558788 515148 558794 515160
rect 559374 515148 559380 515160
rect 558788 515120 559380 515148
rect 558788 515108 558794 515120
rect 559374 515108 559380 515120
rect 559432 515108 559438 515160
rect 301774 513748 301780 513800
rect 301832 513788 301838 513800
rect 301832 513760 303292 513788
rect 301832 513748 301838 513760
rect 303264 513720 303292 513760
rect 306098 513720 306104 513732
rect 303264 513692 306104 513720
rect 306098 513680 306104 513692
rect 306156 513680 306162 513732
rect 314286 512252 314292 512304
rect 314344 512292 314350 512304
rect 314562 512292 314568 512304
rect 314344 512264 314568 512292
rect 314344 512252 314350 512264
rect 314562 512252 314568 512264
rect 314620 512252 314626 512304
rect 268838 510892 268844 510944
rect 268896 510932 268902 510944
rect 276382 510932 276388 510944
rect 268896 510904 276388 510932
rect 268896 510892 268902 510904
rect 276382 510892 276388 510904
rect 276440 510892 276446 510944
rect 306190 509668 306196 509720
rect 306248 509708 306254 509720
rect 307570 509708 307576 509720
rect 306248 509680 307576 509708
rect 306248 509668 306254 509680
rect 307570 509668 307576 509680
rect 307628 509708 307634 509720
rect 315482 509708 315488 509720
rect 307628 509680 315488 509708
rect 307628 509668 307634 509680
rect 315482 509668 315488 509680
rect 315540 509668 315546 509720
rect 314286 504880 314292 504892
rect 314247 504852 314292 504880
rect 314286 504840 314292 504852
rect 314344 504840 314350 504892
rect 314289 494615 314347 494621
rect 314289 494581 314301 494615
rect 314335 494612 314347 494615
rect 314378 494612 314384 494624
rect 314335 494584 314384 494612
rect 314335 494581 314347 494584
rect 314289 494575 314347 494581
rect 314378 494572 314384 494584
rect 314436 494572 314442 494624
rect 314286 484276 314292 484288
rect 314247 484248 314292 484276
rect 314286 484236 314292 484248
rect 314344 484236 314350 484288
rect 314289 474011 314347 474017
rect 314289 473977 314301 474011
rect 314335 474008 314347 474011
rect 314378 474008 314384 474020
rect 314335 473980 314384 474008
rect 314335 473977 314347 473980
rect 314289 473971 314347 473977
rect 314378 473968 314384 473980
rect 314436 473968 314442 474020
rect 270034 472540 270040 472592
rect 270092 472580 270098 472592
rect 315482 472580 315488 472592
rect 270092 472552 315488 472580
rect 270092 472540 270098 472552
rect 315482 472540 315488 472552
rect 315540 472540 315546 472592
rect 314286 463672 314292 463684
rect 314247 463644 314292 463672
rect 314286 463632 314292 463644
rect 314344 463632 314350 463684
rect 314289 453407 314347 453413
rect 314289 453373 314301 453407
rect 314335 453404 314347 453407
rect 314378 453404 314384 453416
rect 314335 453376 314384 453404
rect 314335 453373 314347 453376
rect 314289 453367 314347 453373
rect 314378 453364 314384 453376
rect 314436 453364 314442 453416
rect 269298 440104 269304 440156
rect 269356 440144 269362 440156
rect 286226 440144 286232 440156
rect 269356 440116 286232 440144
rect 269356 440104 269362 440116
rect 286226 440104 286232 440116
rect 286284 440104 286290 440156
rect 314286 435752 314292 435804
rect 314344 435752 314350 435804
rect 314304 435724 314332 435752
rect 314378 435724 314384 435736
rect 314304 435696 314384 435724
rect 314378 435684 314384 435696
rect 314436 435684 314442 435736
rect 314378 432732 314384 432744
rect 314339 432704 314384 432732
rect 314378 432692 314384 432704
rect 314436 432692 314442 432744
rect 558822 432488 558828 432540
rect 558880 432528 558886 432540
rect 560754 432528 560760 432540
rect 558880 432500 560760 432528
rect 558880 432488 558886 432500
rect 560754 432488 560760 432500
rect 560812 432488 560818 432540
rect 314378 425388 314384 425400
rect 314339 425360 314384 425388
rect 314378 425348 314384 425360
rect 314436 425348 314442 425400
rect 314286 412156 314292 412208
rect 314344 412196 314350 412208
rect 314470 412196 314476 412208
rect 314344 412168 314476 412196
rect 314344 412156 314350 412168
rect 314470 412156 314476 412168
rect 314528 412156 314534 412208
rect 269298 404812 269304 404864
rect 269356 404852 269362 404864
rect 303890 404852 303896 404864
rect 269356 404824 303896 404852
rect 269356 404812 269362 404824
rect 303890 404812 303896 404824
rect 303948 404812 303954 404864
rect 314194 401888 314200 401940
rect 314252 401928 314258 401940
rect 316218 401928 316224 401940
rect 314252 401900 316224 401928
rect 314252 401888 314258 401900
rect 316218 401888 316224 401900
rect 316276 401888 316282 401940
rect 314378 394544 314384 394596
rect 314436 394544 314442 394596
rect 314396 394460 314424 394544
rect 314378 394408 314384 394460
rect 314436 394408 314442 394460
rect 558730 391552 558736 391604
rect 558788 391592 558794 391604
rect 578786 391592 578792 391604
rect 558788 391564 578792 391592
rect 558788 391552 558794 391564
rect 578786 391552 578792 391564
rect 578844 391552 578850 391604
rect 24946 386316 24952 386368
rect 25004 386356 25010 386368
rect 313734 386356 313740 386368
rect 25004 386328 313740 386356
rect 25004 386316 25010 386328
rect 313734 386316 313740 386328
rect 313792 386356 313798 386368
rect 314194 386356 314200 386368
rect 313792 386328 314200 386356
rect 313792 386316 313798 386328
rect 314194 386316 314200 386328
rect 314252 386316 314258 386368
rect 286226 386248 286232 386300
rect 286284 386288 286290 386300
rect 558822 386288 558828 386300
rect 286284 386260 558828 386288
rect 286284 386248 286290 386260
rect 558822 386248 558828 386260
rect 558880 386248 558886 386300
rect 286226 385704 286232 385756
rect 286284 385744 286290 385756
rect 286686 385744 286692 385756
rect 286284 385716 286692 385744
rect 286284 385704 286290 385716
rect 286686 385704 286692 385716
rect 286744 385704 286750 385756
rect 87690 382644 87696 382696
rect 87748 382684 87754 382696
rect 273898 382684 273904 382696
rect 87748 382656 273904 382684
rect 87748 382644 87754 382656
rect 273898 382644 273904 382656
rect 273956 382644 273962 382696
rect 232130 382576 232136 382628
rect 232188 382616 232194 382628
rect 297266 382616 297272 382628
rect 232188 382588 297272 382616
rect 232188 382576 232194 382588
rect 297266 382576 297272 382588
rect 297324 382576 297330 382628
rect 256050 382508 256056 382560
rect 256108 382548 256114 382560
rect 272334 382548 272340 382560
rect 256108 382520 272340 382548
rect 256108 382508 256114 382520
rect 272334 382508 272340 382520
rect 272392 382508 272398 382560
rect 208026 382372 208032 382424
rect 208084 382412 208090 382424
rect 278222 382412 278228 382424
rect 208084 382384 278228 382412
rect 208084 382372 208090 382384
rect 278222 382372 278228 382384
rect 278280 382412 278286 382424
rect 279602 382412 279608 382424
rect 278280 382384 279608 382412
rect 278280 382372 278286 382384
rect 279602 382372 279608 382384
rect 279660 382372 279666 382424
rect 300946 382372 300952 382424
rect 301004 382412 301010 382424
rect 331490 382412 331496 382424
rect 301004 382384 331496 382412
rect 301004 382372 301010 382384
rect 331490 382372 331496 382384
rect 331548 382372 331554 382424
rect 270126 382304 270132 382356
rect 270184 382344 270190 382356
rect 355594 382344 355600 382356
rect 270184 382316 355600 382344
rect 270184 382304 270190 382316
rect 355594 382304 355600 382316
rect 355652 382304 355658 382356
rect 183922 382236 183928 382288
rect 183980 382276 183986 382288
rect 313642 382276 313648 382288
rect 183980 382248 313648 382276
rect 183980 382236 183986 382248
rect 313642 382236 313648 382248
rect 313700 382276 313706 382288
rect 314930 382276 314936 382288
rect 313700 382248 314936 382276
rect 313700 382236 313706 382248
rect 314930 382236 314936 382248
rect 314988 382236 314994 382288
rect 111794 382168 111800 382220
rect 111852 382208 111858 382220
rect 279694 382208 279700 382220
rect 111852 382180 279700 382208
rect 111852 382168 111858 382180
rect 279694 382168 279700 382180
rect 279752 382208 279758 382220
rect 403618 382208 403624 382220
rect 279752 382180 403624 382208
rect 279752 382168 279758 382180
rect 403618 382168 403624 382180
rect 403676 382168 403682 382220
rect 135898 382100 135904 382152
rect 135956 382140 135962 382152
rect 313826 382140 313832 382152
rect 135956 382112 313832 382140
rect 135956 382100 135962 382112
rect 313826 382100 313832 382112
rect 313884 382140 313890 382152
rect 427722 382140 427728 382152
rect 313884 382112 427728 382140
rect 313884 382100 313890 382112
rect 427722 382100 427728 382112
rect 427780 382100 427786 382152
rect 63770 382032 63776 382084
rect 63828 382072 63834 382084
rect 270126 382072 270132 382084
rect 63828 382044 270132 382072
rect 63828 382032 63834 382044
rect 270126 382032 270132 382044
rect 270184 382032 270190 382084
rect 279602 382032 279608 382084
rect 279660 382072 279666 382084
rect 499850 382072 499856 382084
rect 279660 382044 499856 382072
rect 279660 382032 279666 382044
rect 499850 382032 499856 382044
rect 499908 382032 499914 382084
rect 39666 381964 39672 382016
rect 39724 382004 39730 382016
rect 300946 382004 300952 382016
rect 39724 381976 300952 382004
rect 39724 381964 39730 381976
rect 300946 381964 300952 381976
rect 301004 381964 301010 382016
rect 314930 381964 314936 382016
rect 314988 382004 314994 382016
rect 475930 382004 475936 382016
rect 314988 381976 475936 382004
rect 314988 381964 314994 381976
rect 475930 381964 475936 381976
rect 475988 381964 475994 382016
rect 314194 373940 314200 373992
rect 314252 373940 314258 373992
rect 314212 373912 314240 373940
rect 314286 373912 314292 373924
rect 314212 373884 314292 373912
rect 314286 373872 314292 373884
rect 314344 373872 314350 373924
rect 314102 360680 314108 360732
rect 314160 360720 314166 360732
rect 314378 360720 314384 360732
rect 314160 360692 314384 360720
rect 314160 360680 314166 360692
rect 314378 360680 314384 360692
rect 314436 360680 314442 360732
rect 273530 359184 273536 359236
rect 273588 359224 273594 359236
rect 278498 359224 278504 359236
rect 273588 359196 278504 359224
rect 273588 359184 273594 359196
rect 278498 359184 278504 359196
rect 278556 359184 278562 359236
rect 299014 358844 299020 358896
rect 299072 358884 299078 358896
rect 300210 358884 300216 358896
rect 299072 358856 300216 358884
rect 299072 358844 299078 358856
rect 300210 358844 300216 358856
rect 300268 358844 300274 358896
rect 305270 358504 305276 358556
rect 305328 358544 305334 358556
rect 558638 358544 558644 358556
rect 305328 358516 558644 358544
rect 305328 358504 305334 358516
rect 558638 358504 558644 358516
rect 558696 358504 558702 358556
rect 284754 358436 284760 358488
rect 284812 358476 284818 358488
rect 294966 358476 294972 358488
rect 284812 358448 294972 358476
rect 284812 358436 284818 358448
rect 294966 358436 294972 358448
rect 295024 358436 295030 358488
rect 303246 358436 303252 358488
rect 303304 358476 303310 358488
rect 579246 358476 579252 358488
rect 303304 358448 579252 358476
rect 303304 358436 303310 358448
rect 579246 358436 579252 358448
rect 579304 358436 579310 358488
rect 282638 358368 282644 358420
rect 282696 358408 282702 358420
rect 579430 358408 579436 358420
rect 282696 358380 579436 358408
rect 282696 358368 282702 358380
rect 579430 358368 579436 358380
rect 579488 358368 579494 358420
rect 24946 357892 24952 357944
rect 25004 357932 25010 357944
rect 311342 357932 311348 357944
rect 25004 357904 311348 357932
rect 25004 357892 25010 357904
rect 311342 357892 311348 357904
rect 311400 357892 311406 357944
rect 273162 357824 273168 357876
rect 273220 357864 273226 357876
rect 296990 357864 296996 357876
rect 273220 357836 296996 357864
rect 273220 357824 273226 357836
rect 296990 357824 296996 357836
rect 297048 357824 297054 357876
rect 147122 357756 147128 357808
rect 147180 357796 147186 357808
rect 284662 357796 284668 357808
rect 147180 357768 284668 357796
rect 147180 357756 147186 357768
rect 284662 357756 284668 357768
rect 284720 357756 284726 357808
rect 309594 354832 309600 354884
rect 309652 354872 309658 354884
rect 312722 354872 312728 354884
rect 309652 354844 312728 354872
rect 309652 354832 309658 354844
rect 312722 354832 312728 354844
rect 312780 354832 312786 354884
rect 3878 354084 3884 354136
rect 3936 354124 3942 354136
rect 311526 354124 311532 354136
rect 3936 354096 311532 354124
rect 3936 354084 3942 354096
rect 311526 354084 311532 354096
rect 311584 354084 311590 354136
rect 270310 354016 270316 354068
rect 270368 354056 270374 354068
rect 579338 354056 579344 354068
rect 270368 354028 579344 354056
rect 270368 354016 270374 354028
rect 579338 354016 579344 354028
rect 579396 354016 579402 354068
rect 3786 353948 3792 354000
rect 3844 353988 3850 354000
rect 313550 353988 313556 354000
rect 3844 353960 313556 353988
rect 3844 353948 3850 353960
rect 313550 353948 313556 353960
rect 313608 353948 313614 354000
rect 314378 353376 314384 353388
rect 314304 353348 314384 353376
rect 314304 353252 314332 353348
rect 314378 353336 314384 353348
rect 314436 353336 314442 353388
rect 269850 353200 269856 353252
rect 269908 353240 269914 353252
rect 270126 353240 270132 353252
rect 269908 353212 270132 353240
rect 269908 353200 269914 353212
rect 270126 353200 270132 353212
rect 270184 353200 270190 353252
rect 314286 353200 314292 353252
rect 314344 353200 314350 353252
rect 269850 350316 269856 350328
rect 269811 350288 269856 350316
rect 269850 350276 269856 350288
rect 269908 350276 269914 350328
rect 272889 343043 272947 343049
rect 272889 343009 272901 343043
rect 272935 343040 272947 343043
rect 272978 343040 272984 343052
rect 272935 343012 272984 343040
rect 272935 343009 272947 343012
rect 272889 343003 272947 343009
rect 272978 343000 272984 343012
rect 273036 343000 273042 343052
rect 314102 343000 314108 343052
rect 314160 343040 314166 343052
rect 314286 343040 314292 343052
rect 314160 343012 314292 343040
rect 314160 343000 314166 343012
rect 314286 343000 314292 343012
rect 314344 343000 314350 343052
rect 272610 342388 272616 342440
rect 272668 342428 272674 342440
rect 272978 342428 272984 342440
rect 272668 342400 272984 342428
rect 272668 342388 272674 342400
rect 272978 342388 272984 342400
rect 273036 342388 273042 342440
rect 269853 340051 269911 340057
rect 269853 340017 269865 340051
rect 269899 340048 269911 340051
rect 269942 340048 269948 340060
rect 269899 340020 269948 340048
rect 269899 340017 269911 340020
rect 269853 340011 269911 340017
rect 269942 340008 269948 340020
rect 270000 340008 270006 340060
rect 272886 340048 272892 340060
rect 272847 340020 272892 340048
rect 272886 340008 272892 340020
rect 272944 340008 272950 340060
rect 268562 339940 268568 339992
rect 268620 339980 268626 339992
rect 269666 339980 269672 339992
rect 268620 339952 269672 339980
rect 268620 339940 268626 339952
rect 269666 339940 269672 339952
rect 269724 339940 269730 339992
rect 314930 334092 314936 334144
rect 314988 334132 314994 334144
rect 558546 334132 558552 334144
rect 314988 334104 558552 334132
rect 314988 334092 314994 334104
rect 558546 334092 558552 334104
rect 558604 334092 558610 334144
rect 268562 329740 268568 329792
rect 268620 329780 268626 329792
rect 269390 329780 269396 329792
rect 268620 329752 269396 329780
rect 268620 329740 268626 329752
rect 269390 329740 269396 329752
rect 269448 329740 269454 329792
rect 3602 313488 3608 313540
rect 3660 313528 3666 313540
rect 308582 313528 308588 313540
rect 3660 313500 308588 313528
rect 3660 313488 3666 313500
rect 308582 313488 308588 313500
rect 308640 313488 308646 313540
rect 3694 313420 3700 313472
rect 3752 313460 3758 313472
rect 285950 313460 285956 313472
rect 3752 313432 285956 313460
rect 3752 313420 3758 313432
rect 285950 313420 285956 313432
rect 286008 313420 286014 313472
rect 292206 313420 292212 313472
rect 292264 313460 292270 313472
rect 579154 313460 579160 313472
rect 292264 313432 579160 313460
rect 292264 313420 292270 313432
rect 579154 313420 579160 313432
rect 579212 313420 579218 313472
rect 24854 313352 24860 313404
rect 24912 313392 24918 313404
rect 273622 313392 273628 313404
rect 24912 313364 273628 313392
rect 24912 313352 24918 313364
rect 273622 313352 273628 313364
rect 273680 313352 273686 313404
rect 287974 313352 287980 313404
rect 288032 313392 288038 313404
rect 558730 313392 558736 313404
rect 288032 313364 558736 313392
rect 288032 313352 288038 313364
rect 558730 313352 558736 313364
rect 558788 313352 558794 313404
rect 122098 312876 122104 312928
rect 122156 312916 122162 312928
rect 289998 312916 290004 312928
rect 122156 312888 290004 312916
rect 122156 312876 122162 312888
rect 289998 312876 290004 312888
rect 290056 312876 290062 312928
rect 98546 312808 98552 312860
rect 98604 312848 98610 312860
rect 300302 312848 300308 312860
rect 98604 312820 300308 312848
rect 98604 312808 98610 312820
rect 300302 312808 300308 312820
rect 300360 312808 300366 312860
rect 24854 312740 24860 312792
rect 24912 312780 24918 312792
rect 302510 312780 302516 312792
rect 24912 312752 302516 312780
rect 24912 312740 24918 312752
rect 302510 312740 302516 312752
rect 302568 312740 302574 312792
rect 270034 312128 270040 312180
rect 270092 312128 270098 312180
rect 270052 312044 270080 312128
rect 270034 311992 270040 312044
rect 270092 311992 270098 312044
rect 270034 309108 270040 309120
rect 269995 309080 270040 309108
rect 270034 309068 270040 309080
rect 270092 309068 270098 309120
rect 269850 297372 269856 297424
rect 269908 297412 269914 297424
rect 270037 297415 270095 297421
rect 270037 297412 270049 297415
rect 269908 297384 270049 297412
rect 269908 297372 269914 297384
rect 270037 297381 270049 297384
rect 270083 297381 270095 297415
rect 270037 297375 270095 297381
rect 269850 293332 269856 293344
rect 269811 293304 269856 293332
rect 269850 293292 269856 293304
rect 269908 293292 269914 293344
rect 269853 287079 269911 287085
rect 269853 287045 269865 287079
rect 269899 287076 269911 287079
rect 269942 287076 269948 287088
rect 269899 287048 269948 287076
rect 269899 287045 269911 287048
rect 269853 287039 269911 287045
rect 269942 287036 269948 287048
rect 270000 287036 270006 287088
rect 97994 276700 98000 276752
rect 98052 276740 98058 276752
rect 98546 276740 98552 276752
rect 98052 276712 98552 276740
rect 98052 276700 98058 276712
rect 98546 276700 98552 276712
rect 98604 276700 98610 276752
rect 278133 276675 278191 276681
rect 278133 276641 278145 276675
rect 278179 276641 278191 276675
rect 278133 276635 278191 276641
rect 278148 276604 278176 276635
rect 288529 276607 288587 276613
rect 288529 276604 288541 276607
rect 204640 276576 214880 276604
rect 278148 276576 288541 276604
rect 188433 276539 188491 276545
rect 188433 276505 188445 276539
rect 188479 276536 188491 276539
rect 188479 276508 200988 276536
rect 188479 276505 188491 276508
rect 188433 276499 188491 276505
rect 200960 276468 200988 276508
rect 204640 276468 204668 276576
rect 214852 276536 214880 276576
rect 288529 276573 288541 276576
rect 288575 276573 288587 276607
rect 288529 276567 288587 276573
rect 214852 276508 214972 276536
rect 214944 276477 214972 276508
rect 200960 276440 204668 276468
rect 214929 276471 214987 276477
rect 214929 276437 214941 276471
rect 214975 276437 214987 276471
rect 214929 276431 214987 276437
rect 225141 276471 225199 276477
rect 225141 276437 225153 276471
rect 225187 276468 225199 276471
rect 257617 276471 257675 276477
rect 225187 276440 229692 276468
rect 225187 276437 225199 276440
rect 225141 276431 225199 276437
rect 188433 276403 188491 276409
rect 188433 276400 188445 276403
rect 188356 276372 188445 276400
rect 146202 276292 146208 276344
rect 146260 276332 146266 276344
rect 147122 276332 147128 276344
rect 146260 276304 147128 276332
rect 146260 276292 146266 276304
rect 147122 276292 147128 276304
rect 147180 276292 147186 276344
rect 188356 276332 188384 276372
rect 188433 276369 188445 276372
rect 188479 276369 188491 276403
rect 229664 276400 229692 276440
rect 237024 276440 247264 276468
rect 237024 276400 237052 276440
rect 229664 276372 237052 276400
rect 188433 276363 188491 276369
rect 178144 276304 188384 276332
rect 195793 276335 195851 276341
rect 177301 276267 177359 276273
rect 177301 276233 177313 276267
rect 177347 276264 177359 276267
rect 178144 276264 178172 276304
rect 195793 276301 195805 276335
rect 195839 276332 195851 276335
rect 204625 276335 204683 276341
rect 204625 276332 204637 276335
rect 195839 276304 204637 276332
rect 195839 276301 195851 276304
rect 195793 276295 195851 276301
rect 204625 276301 204637 276304
rect 204671 276301 204683 276335
rect 204625 276295 204683 276301
rect 177347 276236 178172 276264
rect 214929 276267 214987 276273
rect 177347 276233 177359 276236
rect 177301 276227 177359 276233
rect 214929 276233 214941 276267
rect 214975 276264 214987 276267
rect 225141 276267 225199 276273
rect 225141 276264 225153 276267
rect 214975 276236 225153 276264
rect 214975 276233 214987 276236
rect 214929 276227 214987 276233
rect 225141 276233 225153 276236
rect 225187 276233 225199 276267
rect 247236 276264 247264 276440
rect 257617 276437 257629 276471
rect 257663 276468 257675 276471
rect 267829 276471 267887 276477
rect 267829 276468 267841 276471
rect 257663 276440 267841 276468
rect 257663 276437 257675 276440
rect 257617 276431 257675 276437
rect 267829 276437 267841 276440
rect 267875 276437 267887 276471
rect 267829 276431 267887 276437
rect 404817 276471 404875 276477
rect 404817 276437 404829 276471
rect 404863 276468 404875 276471
rect 453393 276471 453451 276477
rect 453393 276468 453405 276471
rect 404863 276440 425468 276468
rect 404863 276437 404875 276440
rect 404817 276431 404875 276437
rect 278133 276403 278191 276409
rect 278133 276400 278145 276403
rect 260484 276372 278145 276400
rect 260484 276332 260512 276372
rect 278133 276369 278145 276372
rect 278179 276369 278191 276403
rect 365714 276400 365720 276412
rect 278133 276363 278191 276369
rect 291396 276372 365720 276400
rect 250272 276304 260512 276332
rect 250272 276264 250300 276304
rect 284018 276292 284024 276344
rect 284076 276332 284082 276344
rect 291396 276332 291424 276372
rect 365714 276360 365720 276372
rect 365772 276360 365778 276412
rect 368017 276403 368075 276409
rect 368017 276369 368029 276403
rect 368063 276400 368075 276403
rect 378229 276403 378287 276409
rect 378229 276400 378241 276403
rect 368063 276372 378241 276400
rect 368063 276369 368075 276372
rect 368017 276363 368075 276369
rect 378229 276369 378241 276372
rect 378275 276369 378287 276403
rect 378229 276363 378287 276369
rect 388625 276403 388683 276409
rect 388625 276369 388637 276403
rect 388671 276400 388683 276403
rect 394513 276403 394571 276409
rect 394513 276400 394525 276403
rect 388671 276372 394525 276400
rect 388671 276369 388683 276372
rect 388625 276363 388683 276369
rect 394513 276369 394525 276372
rect 394559 276369 394571 276403
rect 425440 276400 425468 276440
rect 445956 276440 453405 276468
rect 445956 276400 445984 276440
rect 453393 276437 453405 276440
rect 453439 276437 453451 276471
rect 453393 276431 453451 276437
rect 425440 276372 432828 276400
rect 394513 276363 394571 276369
rect 284076 276304 291424 276332
rect 284076 276292 284082 276304
rect 294322 276292 294328 276344
rect 294380 276332 294386 276344
rect 413922 276332 413928 276344
rect 294380 276304 413928 276332
rect 294380 276292 294386 276304
rect 413922 276292 413928 276304
rect 413980 276292 413986 276344
rect 432800 276332 432828 276372
rect 443012 276372 445984 276400
rect 435637 276335 435695 276341
rect 435637 276332 435649 276335
rect 432800 276304 435649 276332
rect 435637 276301 435649 276304
rect 435683 276301 435695 276335
rect 435637 276295 435695 276301
rect 435729 276335 435787 276341
rect 435729 276301 435741 276335
rect 435775 276332 435787 276335
rect 443012 276332 443040 276372
rect 435775 276304 443040 276332
rect 453393 276335 453451 276341
rect 435775 276301 435787 276304
rect 435729 276295 435787 276301
rect 453393 276301 453405 276335
rect 453439 276332 453451 276335
rect 461946 276332 461952 276344
rect 453439 276304 461952 276332
rect 453439 276301 453451 276304
rect 453393 276295 453451 276301
rect 461946 276292 461952 276304
rect 462004 276292 462010 276344
rect 247236 276236 250300 276264
rect 394513 276267 394571 276273
rect 225141 276227 225199 276233
rect 394513 276233 394525 276267
rect 394559 276264 394571 276267
rect 394559 276236 404768 276264
rect 394559 276233 394571 276236
rect 394513 276227 394571 276233
rect 73890 276156 73896 276208
rect 73948 276196 73954 276208
rect 195793 276199 195851 276205
rect 195793 276196 195805 276199
rect 73948 276168 195805 276196
rect 73948 276156 73954 276168
rect 195793 276165 195805 276168
rect 195839 276165 195851 276199
rect 195793 276159 195851 276165
rect 209685 276199 209743 276205
rect 209685 276165 209697 276199
rect 209731 276196 209743 276199
rect 237006 276196 237012 276208
rect 209731 276168 237012 276196
rect 209731 276165 209743 276168
rect 209685 276159 209743 276165
rect 237006 276156 237012 276168
rect 237064 276156 237070 276208
rect 247218 276156 247224 276208
rect 247276 276196 247282 276208
rect 257617 276199 257675 276205
rect 257617 276196 257629 276199
rect 247276 276168 257629 276196
rect 247276 276156 247282 276168
rect 257617 276165 257629 276168
rect 257663 276165 257675 276199
rect 257617 276159 257675 276165
rect 267829 276199 267887 276205
rect 267829 276165 267841 276199
rect 267875 276196 267887 276199
rect 284018 276196 284024 276208
rect 267875 276168 284024 276196
rect 267875 276165 267887 276168
rect 267829 276159 267887 276165
rect 284018 276156 284024 276168
rect 284076 276156 284082 276208
rect 288529 276199 288587 276205
rect 288529 276165 288541 276199
rect 288575 276196 288587 276199
rect 298002 276196 298008 276208
rect 288575 276168 298008 276196
rect 288575 276165 288587 276168
rect 288529 276159 288587 276165
rect 298002 276156 298008 276168
rect 298060 276196 298066 276208
rect 306193 276199 306251 276205
rect 306193 276196 306205 276199
rect 298060 276168 306205 276196
rect 298060 276156 298066 276168
rect 306193 276165 306205 276168
rect 306239 276165 306251 276199
rect 306193 276159 306251 276165
rect 316405 276199 316463 276205
rect 316405 276165 316417 276199
rect 316451 276196 316463 276199
rect 326801 276199 326859 276205
rect 326801 276196 326813 276199
rect 316451 276168 326813 276196
rect 316451 276165 316463 276168
rect 316405 276159 316463 276165
rect 326801 276165 326813 276168
rect 326847 276165 326859 276199
rect 326801 276159 326859 276165
rect 337013 276199 337071 276205
rect 337013 276165 337025 276199
rect 337059 276196 337071 276199
rect 347409 276199 347467 276205
rect 347409 276196 347421 276199
rect 337059 276168 347421 276196
rect 337059 276165 337071 276168
rect 337013 276159 337071 276165
rect 347409 276165 347421 276168
rect 347455 276165 347467 276199
rect 347409 276159 347467 276165
rect 357621 276199 357679 276205
rect 357621 276165 357633 276199
rect 357667 276196 357679 276199
rect 368017 276199 368075 276205
rect 368017 276196 368029 276199
rect 357667 276168 368029 276196
rect 357667 276165 357679 276168
rect 357621 276159 357679 276165
rect 368017 276165 368029 276168
rect 368063 276165 368075 276199
rect 368017 276159 368075 276165
rect 378229 276199 378287 276205
rect 378229 276165 378241 276199
rect 378275 276196 378287 276199
rect 388625 276199 388683 276205
rect 388625 276196 388637 276199
rect 378275 276168 388637 276196
rect 378275 276165 378287 276168
rect 378229 276159 378287 276165
rect 388625 276165 388637 276168
rect 388671 276165 388683 276199
rect 404740 276196 404768 276236
rect 404817 276199 404875 276205
rect 404817 276196 404829 276199
rect 404740 276168 404829 276196
rect 388625 276159 388683 276165
rect 404817 276165 404829 276168
rect 404863 276165 404875 276199
rect 404817 276159 404875 276165
rect 170122 276088 170128 276140
rect 170180 276128 170186 276140
rect 177301 276131 177359 276137
rect 177301 276128 177313 276131
rect 170180 276100 177313 276128
rect 170180 276088 170186 276100
rect 177301 276097 177313 276100
rect 177347 276097 177359 276131
rect 177301 276091 177359 276097
rect 194226 276088 194232 276140
rect 194284 276128 194290 276140
rect 270402 276128 270408 276140
rect 194284 276100 270408 276128
rect 194284 276088 194290 276100
rect 270402 276088 270408 276100
rect 270460 276128 270466 276140
rect 486050 276128 486056 276140
rect 270460 276100 486056 276128
rect 270460 276088 270466 276100
rect 486050 276088 486056 276100
rect 486108 276088 486114 276140
rect 204625 276063 204683 276069
rect 204625 276029 204637 276063
rect 204671 276060 204683 276063
rect 209685 276063 209743 276069
rect 209685 276060 209697 276063
rect 204671 276032 209697 276060
rect 204671 276029 204683 276032
rect 204625 276023 204683 276029
rect 209685 276029 209697 276032
rect 209731 276029 209743 276063
rect 209685 276023 209743 276029
rect 218330 276020 218336 276072
rect 218388 276060 218394 276072
rect 270218 276060 270224 276072
rect 218388 276032 270224 276060
rect 218388 276020 218394 276032
rect 270218 276020 270224 276032
rect 270276 276060 270282 276072
rect 510154 276060 510160 276072
rect 270276 276032 510160 276060
rect 270276 276020 270282 276032
rect 510154 276020 510160 276032
rect 510212 276020 510218 276072
rect 49970 275952 49976 276004
rect 50028 275992 50034 276004
rect 306834 275992 306840 276004
rect 50028 275964 306840 275992
rect 50028 275952 50034 275964
rect 306834 275952 306840 275964
rect 306892 275992 306898 276004
rect 341794 275992 341800 276004
rect 306892 275964 341800 275992
rect 306892 275952 306898 275964
rect 341794 275952 341800 275964
rect 341852 275952 341858 276004
rect 347409 275995 347467 276001
rect 347409 275961 347421 275995
rect 347455 275992 347467 275995
rect 357621 275995 357679 276001
rect 357621 275992 357633 275995
rect 347455 275964 357633 275992
rect 347455 275961 347467 275964
rect 347409 275955 347467 275961
rect 357621 275961 357633 275964
rect 357667 275961 357679 275995
rect 357621 275955 357679 275961
rect 306193 275927 306251 275933
rect 306193 275893 306205 275927
rect 306239 275924 306251 275927
rect 316405 275927 316463 275933
rect 316405 275924 316417 275927
rect 306239 275896 316417 275924
rect 306239 275893 306251 275896
rect 306193 275887 306251 275893
rect 316405 275893 316417 275896
rect 316451 275893 316463 275927
rect 316405 275887 316463 275893
rect 326801 275927 326859 275933
rect 326801 275893 326813 275927
rect 326847 275924 326859 275927
rect 337013 275927 337071 275933
rect 337013 275924 337025 275927
rect 326847 275896 337025 275924
rect 326847 275893 326859 275896
rect 326801 275887 326859 275893
rect 337013 275893 337025 275896
rect 337059 275893 337071 275927
rect 337013 275887 337071 275893
rect 242434 275340 242440 275392
rect 242492 275380 242498 275392
rect 293586 275380 293592 275392
rect 242492 275352 293592 275380
rect 242492 275340 242498 275352
rect 293586 275340 293592 275352
rect 293644 275380 293650 275392
rect 534258 275380 534264 275392
rect 293644 275352 534264 275380
rect 293644 275340 293650 275352
rect 534258 275340 534264 275352
rect 534316 275340 534322 275392
rect 266354 275272 266360 275324
rect 266412 275312 266418 275324
rect 289814 275312 289820 275324
rect 266412 275284 289820 275312
rect 266412 275272 266418 275284
rect 289814 275272 289820 275284
rect 289872 275312 289878 275324
rect 558178 275312 558184 275324
rect 289872 275284 558184 275312
rect 289872 275272 289878 275284
rect 558178 275272 558184 275284
rect 558236 275272 558242 275324
rect 27246 272348 27252 272400
rect 27304 272388 27310 272400
rect 276658 272388 276664 272400
rect 27304 272360 276664 272388
rect 27304 272348 27310 272360
rect 276658 272348 276664 272360
rect 276716 272348 276722 272400
rect 314378 272348 314384 272400
rect 314436 272388 314442 272400
rect 560846 272388 560852 272400
rect 314436 272360 560852 272388
rect 314436 272348 314442 272360
rect 560846 272348 560852 272360
rect 560904 272348 560910 272400
rect 24762 272076 24768 272128
rect 24820 272116 24826 272128
rect 306834 272116 306840 272128
rect 24820 272088 306840 272116
rect 24820 272076 24826 272088
rect 306834 272076 306840 272088
rect 306892 272076 306898 272128
rect 276566 272008 276572 272060
rect 276624 272048 276630 272060
rect 558546 272048 558552 272060
rect 276624 272020 558552 272048
rect 276624 272008 276630 272020
rect 558546 272008 558552 272020
rect 558604 272008 558610 272060
rect 24670 271940 24676 271992
rect 24728 271980 24734 271992
rect 313734 271980 313740 271992
rect 24728 271952 313740 271980
rect 24728 271940 24734 271952
rect 313734 271940 313740 271952
rect 313792 271940 313798 271992
rect 275922 271736 275928 271788
rect 275980 271776 275986 271788
rect 276566 271776 276572 271788
rect 275980 271748 276572 271776
rect 275980 271736 275986 271748
rect 276566 271736 276572 271748
rect 276624 271736 276630 271788
rect 313734 270852 313740 270904
rect 313792 270892 313798 270904
rect 314286 270892 314292 270904
rect 313792 270864 314292 270892
rect 313792 270852 313798 270864
rect 314286 270852 314292 270864
rect 314344 270852 314350 270904
rect 276658 270784 276664 270836
rect 276716 270824 276722 270836
rect 315022 270824 315028 270836
rect 276716 270796 315028 270824
rect 276716 270784 276722 270796
rect 315022 270784 315028 270796
rect 315080 270784 315086 270836
rect 268378 238416 268384 238468
rect 268436 238456 268442 238468
rect 314378 238456 314384 238468
rect 268436 238428 314384 238456
rect 268436 238416 268442 238428
rect 314378 238416 314384 238428
rect 314436 238416 314442 238468
rect 270126 236988 270132 237040
rect 270184 237028 270190 237040
rect 270218 237028 270224 237040
rect 270184 237000 270224 237028
rect 270184 236988 270190 237000
rect 270218 236988 270224 237000
rect 270276 236988 270282 237040
rect 270218 226720 270224 226772
rect 270276 226760 270282 226772
rect 270402 226760 270408 226772
rect 270276 226732 270408 226760
rect 270276 226720 270282 226732
rect 270402 226720 270408 226732
rect 270460 226720 270466 226772
rect 270126 216384 270132 216436
rect 270184 216424 270190 216436
rect 270218 216424 270224 216436
rect 270184 216396 270224 216424
rect 270184 216384 270190 216396
rect 270218 216384 270224 216396
rect 270276 216384 270282 216436
rect 558546 206048 558552 206100
rect 558604 206088 558610 206100
rect 558914 206088 558920 206100
rect 558604 206060 558920 206088
rect 558604 206048 558610 206060
rect 558914 206048 558920 206060
rect 558972 206048 558978 206100
rect 268378 202784 268384 202836
rect 268436 202824 268442 202836
rect 275922 202824 275928 202836
rect 268436 202796 275928 202824
rect 268436 202784 268442 202796
rect 275922 202784 275928 202796
rect 275980 202784 275986 202836
rect 306834 200132 306840 200184
rect 306892 200172 306898 200184
rect 315022 200172 315028 200184
rect 306892 200144 315028 200172
rect 306892 200132 306898 200144
rect 315022 200132 315028 200144
rect 315080 200132 315086 200184
rect 270218 195888 270224 195900
rect 270144 195860 270224 195888
rect 270144 195832 270172 195860
rect 270218 195848 270224 195860
rect 270276 195848 270282 195900
rect 270126 195780 270132 195832
rect 270184 195780 270190 195832
rect 270218 185512 270224 185564
rect 270276 185552 270282 185564
rect 270402 185552 270408 185564
rect 270276 185524 270408 185552
rect 270276 185512 270282 185524
rect 270402 185512 270408 185524
rect 270460 185512 270466 185564
rect 269942 175176 269948 175228
rect 270000 175216 270006 175228
rect 270126 175216 270132 175228
rect 270000 175188 270132 175216
rect 270000 175176 270006 175188
rect 270126 175176 270132 175188
rect 270184 175176 270190 175228
rect 270218 164840 270224 164892
rect 270276 164880 270282 164892
rect 270402 164880 270408 164892
rect 270276 164852 270408 164880
rect 270276 164840 270282 164852
rect 270402 164840 270408 164852
rect 270460 164840 270466 164892
rect 312722 164772 312728 164824
rect 312780 164812 312786 164824
rect 315022 164812 315028 164824
rect 312780 164784 315028 164812
rect 312780 164772 312786 164784
rect 315022 164772 315028 164784
rect 315080 164772 315086 164824
rect 270126 157428 270132 157480
rect 270184 157468 270190 157480
rect 270402 157468 270408 157480
rect 270184 157440 270408 157468
rect 270184 157428 270190 157440
rect 270402 157428 270408 157440
rect 270460 157428 270466 157480
rect 270126 152912 270132 152924
rect 270087 152884 270132 152912
rect 270126 152872 270132 152884
rect 270184 152872 270190 152924
rect 270129 144279 270187 144285
rect 270129 144245 270141 144279
rect 270175 144276 270187 144279
rect 270218 144276 270224 144288
rect 270175 144248 270224 144276
rect 270175 144245 270187 144248
rect 270129 144239 270187 144245
rect 270218 144236 270224 144248
rect 270276 144236 270282 144288
rect 270126 131016 270132 131028
rect 270087 130988 270132 131016
rect 270126 130976 270132 130988
rect 270184 130976 270190 131028
rect 267918 130228 267924 130280
rect 267976 130268 267982 130280
rect 286226 130268 286232 130280
rect 267976 130240 286232 130268
rect 267976 130228 267982 130240
rect 286226 130228 286232 130240
rect 286284 130228 286290 130280
rect 270129 120751 270187 120757
rect 270129 120717 270141 120751
rect 270175 120748 270187 120751
rect 270218 120748 270224 120760
rect 270175 120720 270224 120748
rect 270175 120717 270187 120720
rect 270129 120711 270187 120717
rect 270218 120708 270224 120720
rect 270276 120708 270282 120760
rect 558546 119212 558552 119264
rect 558604 119252 558610 119264
rect 559374 119252 559380 119264
rect 558604 119224 559380 119252
rect 558604 119212 558610 119224
rect 559374 119212 559380 119224
rect 559432 119212 559438 119264
rect 270218 116288 270224 116340
rect 270276 116288 270282 116340
rect 270236 116192 270264 116288
rect 270310 116192 270316 116204
rect 270236 116164 270316 116192
rect 270310 116152 270316 116164
rect 270368 116152 270374 116204
rect 286226 114792 286232 114844
rect 286284 114832 286290 114844
rect 286284 114804 287100 114832
rect 286284 114792 286290 114804
rect 287072 114764 287100 114804
rect 289538 114764 289544 114776
rect 287072 114736 289544 114764
rect 289538 114724 289544 114736
rect 289596 114724 289602 114776
rect 289538 111800 289544 111852
rect 289596 111840 289602 111852
rect 292850 111840 292856 111852
rect 289596 111812 292856 111840
rect 289596 111800 289602 111812
rect 292850 111800 292856 111812
rect 292908 111800 292914 111852
rect 292850 109896 292856 109948
rect 292908 109936 292914 109948
rect 294414 109936 294420 109948
rect 292908 109908 294420 109936
rect 292908 109896 292914 109908
rect 294414 109896 294420 109908
rect 294472 109896 294478 109948
rect 294414 108876 294420 108928
rect 294472 108916 294478 108928
rect 297266 108916 297272 108928
rect 294472 108888 297272 108916
rect 294472 108876 294478 108888
rect 297266 108876 297272 108888
rect 297324 108876 297330 108928
rect 270218 101600 270224 101652
rect 270276 101640 270282 101652
rect 270310 101640 270316 101652
rect 270276 101612 270316 101640
rect 270276 101600 270282 101612
rect 270310 101600 270316 101612
rect 270368 101600 270374 101652
rect 297358 97588 297364 97640
rect 297416 97628 297422 97640
rect 298830 97628 298836 97640
rect 297416 97600 298836 97628
rect 297416 97588 297422 97600
rect 298830 97588 298836 97600
rect 298888 97588 298894 97640
rect 267918 94868 267924 94920
rect 267976 94908 267982 94920
rect 303246 94908 303252 94920
rect 267976 94880 303252 94908
rect 267976 94868 267982 94880
rect 303246 94868 303252 94880
rect 303304 94908 303310 94920
rect 303890 94908 303896 94920
rect 303304 94880 303896 94908
rect 303304 94868 303310 94880
rect 303890 94868 303896 94880
rect 303948 94868 303954 94920
rect 314194 92352 314200 92404
rect 314252 92392 314258 92404
rect 315022 92392 315028 92404
rect 314252 92364 315028 92392
rect 314252 92352 314258 92364
rect 315022 92352 315028 92364
rect 315080 92352 315086 92404
rect 270034 91264 270040 91316
rect 270092 91304 270098 91316
rect 270126 91304 270132 91316
rect 270092 91276 270132 91304
rect 270092 91264 270098 91276
rect 270126 91264 270132 91276
rect 270184 91264 270190 91316
rect 298830 89768 298836 89820
rect 298888 89808 298894 89820
rect 298888 89780 300348 89808
rect 298888 89768 298894 89780
rect 300320 89740 300348 89780
rect 301774 89740 301780 89752
rect 300320 89712 301780 89740
rect 301774 89700 301780 89712
rect 301832 89700 301838 89752
rect 301774 86912 301780 86964
rect 301832 86952 301838 86964
rect 301832 86924 304764 86952
rect 301832 86912 301838 86924
rect 304736 86816 304764 86924
rect 308950 86816 308956 86828
rect 304736 86788 308956 86816
rect 308950 86776 308956 86788
rect 309008 86776 309014 86828
rect 308950 84192 308956 84244
rect 309008 84232 309014 84244
rect 312078 84232 312084 84244
rect 309008 84204 312084 84232
rect 309008 84192 309014 84204
rect 312078 84192 312084 84204
rect 312136 84192 312142 84244
rect 269666 82356 269672 82408
rect 269724 82396 269730 82408
rect 269942 82396 269948 82408
rect 269724 82368 269948 82396
rect 269724 82356 269730 82368
rect 269942 82356 269948 82368
rect 270000 82356 270006 82408
rect 312078 80928 312084 80980
rect 312136 80968 312142 80980
rect 316402 80968 316408 80980
rect 312136 80940 316408 80968
rect 312136 80928 312142 80940
rect 316402 80928 316408 80940
rect 316460 80928 316466 80980
rect 24946 75964 24952 76016
rect 25004 76004 25010 76016
rect 314194 76004 314200 76016
rect 25004 75976 314200 76004
rect 25004 75964 25010 75976
rect 314194 75964 314200 75976
rect 314252 75964 314258 76016
rect 316494 75964 316500 76016
rect 316552 76004 316558 76016
rect 558546 76004 558552 76016
rect 316552 75976 558552 76004
rect 316552 75964 316558 75976
rect 558546 75964 558552 75976
rect 558604 75964 558610 76016
rect 303890 75896 303896 75948
rect 303948 75936 303954 75948
rect 560846 75936 560852 75948
rect 303948 75908 560852 75936
rect 303948 75896 303954 75908
rect 560846 75896 560852 75908
rect 560904 75896 560910 75948
rect 256050 72088 256056 72140
rect 256108 72128 256114 72140
rect 269761 72131 269819 72137
rect 269761 72128 269773 72131
rect 256108 72100 269773 72128
rect 256108 72088 256114 72100
rect 269761 72097 269773 72100
rect 269807 72097 269819 72131
rect 269761 72091 269819 72097
rect 270037 72131 270095 72137
rect 270037 72097 270049 72131
rect 270083 72128 270095 72131
rect 279694 72128 279700 72140
rect 270083 72100 279700 72128
rect 270083 72097 270095 72100
rect 270037 72091 270095 72097
rect 279694 72088 279700 72100
rect 279752 72128 279758 72140
rect 548058 72128 548064 72140
rect 279752 72100 548064 72128
rect 279752 72088 279758 72100
rect 548058 72088 548064 72100
rect 548116 72088 548122 72140
rect 39666 72020 39672 72072
rect 39724 72060 39730 72072
rect 300946 72060 300952 72072
rect 39724 72032 300952 72060
rect 39724 72020 39730 72032
rect 300946 72020 300952 72032
rect 301004 72020 301010 72072
rect 313642 72020 313648 72072
rect 313700 72060 313706 72072
rect 475930 72060 475936 72072
rect 313700 72032 475936 72060
rect 313700 72020 313706 72032
rect 475930 72020 475936 72032
rect 475988 72020 475994 72072
rect 87690 71952 87696 72004
rect 87748 71992 87754 72004
rect 281166 71992 281172 72004
rect 87748 71964 281172 71992
rect 87748 71952 87754 71964
rect 281166 71952 281172 71964
rect 281224 71952 281230 72004
rect 296070 71952 296076 72004
rect 296128 71992 296134 72004
rect 296530 71992 296536 72004
rect 296128 71964 296536 71992
rect 296128 71952 296134 71964
rect 296530 71952 296536 71964
rect 296588 71992 296594 72004
rect 523954 71992 523960 72004
rect 296588 71964 523960 71992
rect 296588 71952 296594 71964
rect 523954 71952 523960 71964
rect 524012 71952 524018 72004
rect 160002 71884 160008 71936
rect 160060 71924 160066 71936
rect 273162 71924 273168 71936
rect 160060 71896 273168 71924
rect 160060 71884 160066 71896
rect 273162 71884 273168 71896
rect 273220 71884 273226 71936
rect 273254 71884 273260 71936
rect 273312 71924 273318 71936
rect 273530 71924 273536 71936
rect 273312 71896 273536 71924
rect 273312 71884 273318 71896
rect 273530 71884 273536 71896
rect 273588 71924 273594 71936
rect 499850 71924 499856 71936
rect 273588 71896 499856 71924
rect 273588 71884 273594 71896
rect 499850 71884 499856 71896
rect 499908 71884 499914 71936
rect 135898 71816 135904 71868
rect 135956 71856 135962 71868
rect 313550 71856 313556 71868
rect 135956 71828 313556 71856
rect 135956 71816 135962 71828
rect 313550 71816 313556 71828
rect 313608 71856 313614 71868
rect 427722 71856 427728 71868
rect 313608 71828 427728 71856
rect 313608 71816 313614 71828
rect 427722 71816 427728 71828
rect 427780 71816 427786 71868
rect 111794 71748 111800 71800
rect 111852 71788 111858 71800
rect 276658 71788 276664 71800
rect 111852 71760 276664 71788
rect 111852 71748 111858 71760
rect 276658 71748 276664 71760
rect 276716 71788 276722 71800
rect 403618 71788 403624 71800
rect 276716 71760 403624 71788
rect 276716 71748 276722 71760
rect 403618 71748 403624 71760
rect 403676 71748 403682 71800
rect 183922 71680 183928 71732
rect 183980 71720 183986 71732
rect 313642 71720 313648 71732
rect 183980 71692 313648 71720
rect 183980 71680 183986 71692
rect 313642 71680 313648 71692
rect 313700 71680 313706 71732
rect 208026 71612 208032 71664
rect 208084 71652 208090 71664
rect 273254 71652 273260 71664
rect 208084 71624 273260 71652
rect 208084 71612 208090 71624
rect 273254 71612 273260 71624
rect 273312 71612 273318 71664
rect 281166 71612 281172 71664
rect 281224 71652 281230 71664
rect 379514 71652 379520 71664
rect 281224 71624 379520 71652
rect 281224 71612 281230 71624
rect 379514 71612 379520 71624
rect 379572 71612 379578 71664
rect 63770 71544 63776 71596
rect 63828 71584 63834 71596
rect 269758 71584 269764 71596
rect 63828 71556 269764 71584
rect 63828 71544 63834 71556
rect 269758 71544 269764 71556
rect 269816 71584 269822 71596
rect 355594 71584 355600 71596
rect 269816 71556 355600 71584
rect 269816 71544 269822 71556
rect 355594 71544 355600 71556
rect 355652 71544 355658 71596
rect 232130 71476 232136 71528
rect 232188 71516 232194 71528
rect 296070 71516 296076 71528
rect 232188 71488 296076 71516
rect 232188 71476 232194 71488
rect 296070 71476 296076 71488
rect 296128 71476 296134 71528
rect 300946 71476 300952 71528
rect 301004 71516 301010 71528
rect 331490 71516 331496 71528
rect 301004 71488 331496 71516
rect 301004 71476 301010 71488
rect 331490 71476 331496 71488
rect 331548 71476 331554 71528
rect 270586 3612 270592 3664
rect 270644 3652 270650 3664
rect 583386 3652 583392 3664
rect 270644 3624 583392 3652
rect 270644 3612 270650 3624
rect 583386 3612 583392 3624
rect 583444 3612 583450 3664
<< via1 >>
rect 8024 700612 8076 700664
rect 8208 700612 8260 700664
rect 72976 700612 73028 700664
rect 137836 700612 137888 700664
rect 202788 700612 202840 700664
rect 267648 700612 267700 700664
rect 273812 700612 273864 700664
rect 332508 700612 332560 700664
rect 397460 700612 397512 700664
rect 462320 700612 462372 700664
rect 527180 700612 527232 700664
rect 272984 700068 273036 700120
rect 283840 700068 283892 700120
rect 273076 700000 273128 700052
rect 364984 700000 365036 700052
rect 270684 699932 270736 699984
rect 429844 699932 429896 699984
rect 527180 699932 527232 699984
rect 579896 699932 579948 699984
rect 154120 699864 154172 699916
rect 268568 699864 268620 699916
rect 270776 699864 270828 699916
rect 559656 699864 559708 699916
rect 2964 653488 3016 653540
rect 8024 653488 8076 653540
rect 270500 627104 270552 627156
rect 578792 627104 578844 627156
rect 49608 586440 49660 586492
rect 307576 586440 307628 586492
rect 73528 586372 73580 586424
rect 289452 586372 289504 586424
rect 485780 586440 485832 586492
rect 219348 586304 219400 586356
rect 242072 586304 242124 586356
rect 293592 586304 293644 586356
rect 169760 586236 169812 586288
rect 298652 586236 298704 586288
rect 193864 586100 193916 586152
rect 270408 586100 270460 586152
rect 270592 586100 270644 586152
rect 509884 586100 509936 586152
rect 145840 586032 145892 586084
rect 284760 586032 284812 586084
rect 293592 586032 293644 586084
rect 533988 586032 534040 586084
rect 217968 585964 218020 586016
rect 270592 585964 270644 586016
rect 300216 585964 300268 586016
rect 437756 585964 437808 586016
rect 219348 585896 219400 585948
rect 265992 585896 266044 585948
rect 289176 585896 289228 585948
rect 557908 585896 557960 585948
rect 24860 582428 24912 582480
rect 314384 582428 314436 582480
rect 26516 582360 26568 582412
rect 267096 582360 267148 582412
rect 27252 582292 27304 582344
rect 276664 582292 276716 582344
rect 319444 582292 319496 582344
rect 558736 582292 558788 582344
rect 313464 582224 313516 582276
rect 560852 582224 560904 582276
rect 276664 580660 276716 580712
rect 315396 580660 315448 580712
rect 558552 579980 558604 580032
rect 578792 579980 578844 580032
rect 317972 578484 318024 578536
rect 319444 578484 319496 578536
rect 267096 575492 267148 575544
rect 271880 575492 271932 575544
rect 24952 573996 25004 574048
rect 26516 574064 26568 574116
rect 309140 573996 309192 574048
rect 317972 574064 318024 574116
rect 305368 571820 305420 571872
rect 309140 571820 309192 571872
rect 271880 571208 271932 571260
rect 276572 571072 276624 571124
rect 276572 566652 276624 566704
rect 279240 566652 279292 566704
rect 314108 565224 314160 565276
rect 314384 565224 314436 565276
rect 279240 560056 279292 560108
rect 280344 560056 280396 560108
rect 301688 557812 301740 557864
rect 305368 557880 305420 557932
rect 299572 554344 299624 554396
rect 301688 554344 301740 554396
rect 297364 552032 297416 552084
rect 299572 552032 299624 552084
rect 268292 548972 268344 549024
rect 313464 548972 313516 549024
rect 313464 547612 313516 547664
rect 313924 547612 313976 547664
rect 314200 544824 314252 544876
rect 315856 544824 315908 544876
rect 295892 543736 295944 543788
rect 297364 543736 297416 543788
rect 280344 538704 280396 538756
rect 282184 538704 282236 538756
rect 294420 538024 294472 538076
rect 295892 538024 295944 538076
rect 282184 535032 282236 535084
rect 288532 535032 288584 535084
rect 288532 533944 288584 533996
rect 290004 533944 290056 533996
rect 291384 533672 291436 533724
rect 294420 533672 294472 533724
rect 558644 532856 558696 532908
rect 578792 532856 578844 532908
rect 289268 528436 289320 528488
rect 291384 528436 291436 528488
rect 290004 526940 290056 526992
rect 292764 526940 292816 526992
rect 292764 524016 292816 524068
rect 295524 523948 295576 524000
rect 287060 523200 287112 523252
rect 289268 523200 289320 523252
rect 295524 521024 295576 521076
rect 298468 521024 298520 521076
rect 284116 516672 284168 516724
rect 286968 516672 287020 516724
rect 298468 516672 298520 516724
rect 301780 516672 301832 516724
rect 283288 515176 283340 515228
rect 284116 515176 284168 515228
rect 558736 515108 558788 515160
rect 559380 515108 559432 515160
rect 301780 513748 301832 513800
rect 306104 513680 306156 513732
rect 314292 512252 314344 512304
rect 314568 512252 314620 512304
rect 268844 510892 268896 510944
rect 276388 510892 276440 510944
rect 306196 509668 306248 509720
rect 307576 509668 307628 509720
rect 315488 509668 315540 509720
rect 314292 504883 314344 504892
rect 314292 504849 314301 504883
rect 314301 504849 314335 504883
rect 314335 504849 314344 504883
rect 314292 504840 314344 504849
rect 314384 494572 314436 494624
rect 314292 484279 314344 484288
rect 314292 484245 314301 484279
rect 314301 484245 314335 484279
rect 314335 484245 314344 484279
rect 314292 484236 314344 484245
rect 314384 473968 314436 474020
rect 270040 472540 270092 472592
rect 315488 472540 315540 472592
rect 314292 463675 314344 463684
rect 314292 463641 314301 463675
rect 314301 463641 314335 463675
rect 314335 463641 314344 463675
rect 314292 463632 314344 463641
rect 314384 453364 314436 453416
rect 269304 440104 269356 440156
rect 286232 440104 286284 440156
rect 314292 435752 314344 435804
rect 314384 435684 314436 435736
rect 314384 432735 314436 432744
rect 314384 432701 314393 432735
rect 314393 432701 314427 432735
rect 314427 432701 314436 432735
rect 314384 432692 314436 432701
rect 558828 432488 558880 432540
rect 560760 432488 560812 432540
rect 314384 425391 314436 425400
rect 314384 425357 314393 425391
rect 314393 425357 314427 425391
rect 314427 425357 314436 425391
rect 314384 425348 314436 425357
rect 314292 412156 314344 412208
rect 314476 412156 314528 412208
rect 269304 404812 269356 404864
rect 303896 404812 303948 404864
rect 314200 401888 314252 401940
rect 316224 401888 316276 401940
rect 314384 394544 314436 394596
rect 314384 394408 314436 394460
rect 558736 391552 558788 391604
rect 578792 391552 578844 391604
rect 24952 386316 25004 386368
rect 313740 386316 313792 386368
rect 314200 386316 314252 386368
rect 286232 386248 286284 386300
rect 558828 386248 558880 386300
rect 286232 385704 286284 385756
rect 286692 385704 286744 385756
rect 87696 382644 87748 382696
rect 273904 382644 273956 382696
rect 232136 382576 232188 382628
rect 297272 382576 297324 382628
rect 256056 382508 256108 382560
rect 272340 382508 272392 382560
rect 208032 382372 208084 382424
rect 278228 382372 278280 382424
rect 279608 382372 279660 382424
rect 300952 382372 301004 382424
rect 331496 382372 331548 382424
rect 270132 382304 270184 382356
rect 355600 382304 355652 382356
rect 183928 382236 183980 382288
rect 313648 382236 313700 382288
rect 314936 382236 314988 382288
rect 111800 382168 111852 382220
rect 279700 382168 279752 382220
rect 403624 382168 403676 382220
rect 135904 382100 135956 382152
rect 313832 382100 313884 382152
rect 427728 382100 427780 382152
rect 63776 382032 63828 382084
rect 270132 382032 270184 382084
rect 279608 382032 279660 382084
rect 499856 382032 499908 382084
rect 39672 381964 39724 382016
rect 300952 381964 301004 382016
rect 314936 381964 314988 382016
rect 475936 381964 475988 382016
rect 314200 373940 314252 373992
rect 314292 373872 314344 373924
rect 314108 360680 314160 360732
rect 314384 360680 314436 360732
rect 273536 359184 273588 359236
rect 278504 359184 278556 359236
rect 299020 358844 299072 358896
rect 300216 358844 300268 358896
rect 305276 358504 305328 358556
rect 558644 358504 558696 358556
rect 284760 358436 284812 358488
rect 294972 358436 295024 358488
rect 303252 358436 303304 358488
rect 579252 358436 579304 358488
rect 282644 358368 282696 358420
rect 579436 358368 579488 358420
rect 24952 357892 25004 357944
rect 311348 357892 311400 357944
rect 273168 357824 273220 357876
rect 296996 357824 297048 357876
rect 147128 357756 147180 357808
rect 284668 357756 284720 357808
rect 309600 354832 309652 354884
rect 312728 354832 312780 354884
rect 3884 354084 3936 354136
rect 311532 354084 311584 354136
rect 270316 354016 270368 354068
rect 579344 354016 579396 354068
rect 3792 353948 3844 354000
rect 313556 353948 313608 354000
rect 314384 353336 314436 353388
rect 269856 353200 269908 353252
rect 270132 353200 270184 353252
rect 314292 353200 314344 353252
rect 269856 350319 269908 350328
rect 269856 350285 269865 350319
rect 269865 350285 269899 350319
rect 269899 350285 269908 350319
rect 269856 350276 269908 350285
rect 272984 343000 273036 343052
rect 314108 343000 314160 343052
rect 314292 343000 314344 343052
rect 272616 342388 272668 342440
rect 272984 342388 273036 342440
rect 269948 340008 270000 340060
rect 272892 340051 272944 340060
rect 272892 340017 272901 340051
rect 272901 340017 272935 340051
rect 272935 340017 272944 340051
rect 272892 340008 272944 340017
rect 268568 339940 268620 339992
rect 269672 339940 269724 339992
rect 314936 334092 314988 334144
rect 558552 334092 558604 334144
rect 268568 329740 268620 329792
rect 269396 329740 269448 329792
rect 3608 313488 3660 313540
rect 308588 313488 308640 313540
rect 3700 313420 3752 313472
rect 285956 313420 286008 313472
rect 292212 313420 292264 313472
rect 579160 313420 579212 313472
rect 24860 313352 24912 313404
rect 273628 313352 273680 313404
rect 287980 313352 288032 313404
rect 558736 313352 558788 313404
rect 122104 312876 122156 312928
rect 290004 312876 290056 312928
rect 98552 312808 98604 312860
rect 300308 312808 300360 312860
rect 24860 312740 24912 312792
rect 302516 312740 302568 312792
rect 270040 312128 270092 312180
rect 270040 311992 270092 312044
rect 270040 309111 270092 309120
rect 270040 309077 270049 309111
rect 270049 309077 270083 309111
rect 270083 309077 270092 309111
rect 270040 309068 270092 309077
rect 269856 297372 269908 297424
rect 269856 293335 269908 293344
rect 269856 293301 269865 293335
rect 269865 293301 269899 293335
rect 269899 293301 269908 293335
rect 269856 293292 269908 293301
rect 269948 287036 270000 287088
rect 98000 276700 98052 276752
rect 98552 276700 98604 276752
rect 146208 276292 146260 276344
rect 147128 276292 147180 276344
rect 284024 276292 284076 276344
rect 365720 276360 365772 276412
rect 294328 276292 294380 276344
rect 413928 276292 413980 276344
rect 461952 276292 462004 276344
rect 73896 276156 73948 276208
rect 237012 276156 237064 276208
rect 247224 276156 247276 276208
rect 284024 276156 284076 276208
rect 298008 276156 298060 276208
rect 170128 276088 170180 276140
rect 194232 276088 194284 276140
rect 270408 276088 270460 276140
rect 486056 276088 486108 276140
rect 218336 276020 218388 276072
rect 270224 276020 270276 276072
rect 510160 276020 510212 276072
rect 49976 275952 50028 276004
rect 306840 275952 306892 276004
rect 341800 275952 341852 276004
rect 242440 275340 242492 275392
rect 293592 275340 293644 275392
rect 534264 275340 534316 275392
rect 266360 275272 266412 275324
rect 289820 275272 289872 275324
rect 558184 275272 558236 275324
rect 27252 272348 27304 272400
rect 276664 272348 276716 272400
rect 314384 272348 314436 272400
rect 560852 272348 560904 272400
rect 24768 272076 24820 272128
rect 306840 272076 306892 272128
rect 276572 272008 276624 272060
rect 558552 272008 558604 272060
rect 24676 271940 24728 271992
rect 313740 271940 313792 271992
rect 275928 271736 275980 271788
rect 276572 271736 276624 271788
rect 313740 270852 313792 270904
rect 314292 270852 314344 270904
rect 276664 270784 276716 270836
rect 315028 270784 315080 270836
rect 268384 238416 268436 238468
rect 314384 238416 314436 238468
rect 270132 236988 270184 237040
rect 270224 236988 270276 237040
rect 270224 226720 270276 226772
rect 270408 226720 270460 226772
rect 270132 216384 270184 216436
rect 270224 216384 270276 216436
rect 558552 206048 558604 206100
rect 558920 206048 558972 206100
rect 268384 202784 268436 202836
rect 275928 202784 275980 202836
rect 306840 200132 306892 200184
rect 315028 200132 315080 200184
rect 270224 195848 270276 195900
rect 270132 195780 270184 195832
rect 270224 185512 270276 185564
rect 270408 185512 270460 185564
rect 269948 175176 270000 175228
rect 270132 175176 270184 175228
rect 270224 164840 270276 164892
rect 270408 164840 270460 164892
rect 312728 164772 312780 164824
rect 315028 164772 315080 164824
rect 270132 157428 270184 157480
rect 270408 157428 270460 157480
rect 270132 152915 270184 152924
rect 270132 152881 270141 152915
rect 270141 152881 270175 152915
rect 270175 152881 270184 152915
rect 270132 152872 270184 152881
rect 270224 144236 270276 144288
rect 270132 131019 270184 131028
rect 270132 130985 270141 131019
rect 270141 130985 270175 131019
rect 270175 130985 270184 131019
rect 270132 130976 270184 130985
rect 267924 130228 267976 130280
rect 286232 130228 286284 130280
rect 270224 120708 270276 120760
rect 558552 119212 558604 119264
rect 559380 119212 559432 119264
rect 270224 116288 270276 116340
rect 270316 116152 270368 116204
rect 286232 114792 286284 114844
rect 289544 114724 289596 114776
rect 289544 111800 289596 111852
rect 292856 111800 292908 111852
rect 292856 109896 292908 109948
rect 294420 109896 294472 109948
rect 294420 108876 294472 108928
rect 297272 108876 297324 108928
rect 270224 101600 270276 101652
rect 270316 101600 270368 101652
rect 297364 97588 297416 97640
rect 298836 97588 298888 97640
rect 267924 94868 267976 94920
rect 303252 94868 303304 94920
rect 303896 94868 303948 94920
rect 314200 92352 314252 92404
rect 315028 92352 315080 92404
rect 270040 91264 270092 91316
rect 270132 91264 270184 91316
rect 298836 89768 298888 89820
rect 301780 89700 301832 89752
rect 301780 86912 301832 86964
rect 308956 86776 309008 86828
rect 308956 84192 309008 84244
rect 312084 84192 312136 84244
rect 269672 82356 269724 82408
rect 269948 82356 270000 82408
rect 312084 80928 312136 80980
rect 316408 80928 316460 80980
rect 24952 75964 25004 76016
rect 314200 75964 314252 76016
rect 316500 75964 316552 76016
rect 558552 75964 558604 76016
rect 303896 75896 303948 75948
rect 560852 75896 560904 75948
rect 256056 72088 256108 72140
rect 279700 72088 279752 72140
rect 548064 72088 548116 72140
rect 39672 72020 39724 72072
rect 300952 72020 301004 72072
rect 313648 72020 313700 72072
rect 475936 72020 475988 72072
rect 87696 71952 87748 72004
rect 281172 71952 281224 72004
rect 296076 71952 296128 72004
rect 296536 71952 296588 72004
rect 523960 71952 524012 72004
rect 160008 71884 160060 71936
rect 273168 71884 273220 71936
rect 273260 71884 273312 71936
rect 273536 71884 273588 71936
rect 499856 71884 499908 71936
rect 135904 71816 135956 71868
rect 313556 71816 313608 71868
rect 427728 71816 427780 71868
rect 111800 71748 111852 71800
rect 276664 71748 276716 71800
rect 403624 71748 403676 71800
rect 183928 71680 183980 71732
rect 313648 71680 313700 71732
rect 208032 71612 208084 71664
rect 273260 71612 273312 71664
rect 281172 71612 281224 71664
rect 379520 71612 379572 71664
rect 63776 71544 63828 71596
rect 269764 71544 269816 71596
rect 355600 71544 355652 71596
rect 232136 71476 232188 71528
rect 296076 71476 296128 71528
rect 300952 71476 301004 71528
rect 331496 71476 331548 71528
rect 270592 3612 270644 3664
rect 583392 3612 583444 3664
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 703474 8156 703520
rect 8128 703446 8248 703474
rect 8220 700670 8248 703446
rect 8024 700664 8076 700670
rect 8024 700606 8076 700612
rect 8208 700664 8260 700670
rect 8208 700606 8260 700612
rect 3606 667992 3662 668001
rect 3606 667927 3662 667936
rect 2962 653576 3018 653585
rect 2962 653511 2964 653520
rect 3016 653511 3018 653520
rect 2964 653482 3016 653488
rect 2976 596057 3004 653482
rect 2962 596048 3018 596057
rect 2962 595983 3018 595992
rect 2976 538665 3004 595983
rect 2962 538656 3018 538665
rect 2962 538591 3018 538600
rect 2976 481137 3004 538591
rect 2962 481128 3018 481137
rect 2962 481063 3018 481072
rect 3620 313546 3648 667927
rect 8036 653546 8064 700606
rect 24320 699961 24348 703520
rect 72988 700670 73016 703520
rect 72976 700664 73028 700670
rect 72976 700606 73028 700612
rect 89180 700097 89208 703520
rect 137848 700670 137876 703520
rect 137836 700664 137888 700670
rect 137836 700606 137888 700612
rect 89166 700088 89222 700097
rect 89166 700023 89222 700032
rect 24306 699952 24362 699961
rect 154132 699922 154160 703520
rect 202800 700670 202828 703520
rect 202788 700664 202840 700670
rect 202788 700606 202840 700612
rect 218992 700233 219020 703520
rect 267660 700670 267688 703520
rect 267648 700664 267700 700670
rect 267648 700606 267700 700612
rect 273812 700664 273864 700670
rect 273812 700606 273864 700612
rect 218978 700224 219034 700233
rect 218978 700159 219034 700168
rect 272984 700120 273036 700126
rect 272984 700062 273036 700068
rect 270684 699984 270736 699990
rect 270684 699926 270736 699932
rect 24306 699887 24362 699896
rect 154120 699916 154172 699922
rect 154120 699858 154172 699864
rect 268568 699916 268620 699922
rect 268568 699858 268620 699864
rect 8024 653540 8076 653546
rect 8024 653482 8076 653488
rect 3698 610464 3754 610473
rect 3698 610399 3754 610408
rect 3608 313540 3660 313546
rect 3608 313482 3660 313488
rect 3712 313478 3740 610399
rect 49608 586492 49660 586498
rect 49608 586434 49660 586440
rect 49620 583930 49648 586434
rect 73528 586424 73580 586430
rect 73528 586366 73580 586372
rect 73540 583930 73568 586366
rect 219348 586356 219400 586362
rect 219348 586298 219400 586304
rect 242072 586356 242124 586362
rect 242072 586298 242124 586304
rect 169760 586288 169812 586294
rect 169760 586230 169812 586236
rect 145840 586084 145892 586090
rect 145840 586026 145892 586032
rect 121734 585984 121790 585993
rect 121734 585919 121790 585928
rect 121748 583930 121776 585919
rect 145852 583930 145880 586026
rect 169772 583930 169800 586230
rect 193864 586152 193916 586158
rect 193864 586094 193916 586100
rect 193876 583930 193904 586094
rect 217968 586016 218020 586022
rect 217968 585958 218020 585964
rect 217980 583930 218008 585958
rect 219360 585954 219388 586298
rect 219348 585948 219400 585954
rect 219348 585890 219400 585896
rect 242084 583930 242112 586298
rect 265992 585948 266044 585954
rect 265992 585890 266044 585896
rect 266004 583930 266032 585890
rect 49620 583902 49680 583930
rect 73540 583902 73600 583930
rect 121748 583902 121808 583930
rect 145852 583902 145912 583930
rect 169772 583902 169832 583930
rect 193876 583902 193936 583930
rect 217980 583902 218040 583930
rect 242084 583902 242144 583930
rect 266004 583902 266064 583930
rect 24860 582480 24912 582486
rect 24860 582422 24912 582428
rect 3790 553072 3846 553081
rect 3790 553007 3846 553016
rect 3804 354006 3832 553007
rect 24872 545601 24900 582422
rect 26516 582412 26568 582418
rect 26516 582354 26568 582360
rect 267096 582412 267148 582418
rect 267096 582354 267148 582360
rect 26528 574122 26556 582354
rect 27252 582344 27304 582350
rect 27252 582286 27304 582292
rect 27264 581233 27292 582286
rect 27250 581224 27306 581233
rect 27250 581159 27306 581168
rect 267108 575550 267136 582354
rect 267096 575544 267148 575550
rect 267096 575486 267148 575492
rect 26516 574116 26568 574122
rect 26516 574058 26568 574064
rect 24952 574048 25004 574054
rect 24952 573990 25004 573996
rect 24858 545592 24914 545601
rect 24858 545527 24914 545536
rect 24964 509969 24992 573990
rect 268292 549024 268344 549030
rect 268292 548966 268344 548972
rect 268304 547777 268332 548966
rect 268290 547768 268346 547777
rect 268290 547703 268346 547712
rect 24950 509960 25006 509969
rect 24950 509895 25006 509904
rect 3882 495544 3938 495553
rect 3882 495479 3938 495488
rect 3896 354142 3924 495479
rect 24858 473104 24914 473113
rect 24858 473039 24914 473048
rect 3884 354136 3936 354142
rect 3884 354078 3936 354084
rect 3792 354000 3844 354006
rect 3792 353942 3844 353948
rect 3700 313472 3752 313478
rect 3700 313414 3752 313420
rect 24872 313410 24900 473039
rect 24950 402112 25006 402121
rect 24950 402047 25006 402056
rect 24964 386374 24992 402047
rect 24952 386368 25004 386374
rect 24952 386310 25004 386316
rect 39376 383982 39712 384010
rect 63480 383982 63816 384010
rect 87400 383982 87736 384010
rect 111504 383982 111840 384010
rect 135608 383982 135944 384010
rect 183816 383982 183968 384010
rect 207736 383982 208072 384010
rect 231840 383982 232176 384010
rect 255944 383982 256096 384010
rect 39684 382022 39712 383982
rect 63788 382090 63816 383982
rect 87708 382702 87736 383982
rect 87696 382696 87748 382702
rect 87696 382638 87748 382644
rect 111812 382226 111840 383982
rect 111800 382220 111852 382226
rect 111800 382162 111852 382168
rect 135916 382158 135944 383982
rect 183940 382294 183968 383982
rect 208044 382430 208072 383982
rect 232148 382634 232176 383982
rect 232136 382628 232188 382634
rect 232136 382570 232188 382576
rect 256068 382566 256096 383982
rect 256056 382560 256108 382566
rect 256056 382502 256108 382508
rect 208032 382424 208084 382430
rect 208032 382366 208084 382372
rect 183928 382288 183980 382294
rect 183928 382230 183980 382236
rect 135904 382152 135956 382158
rect 135904 382094 135956 382100
rect 63776 382084 63828 382090
rect 63776 382026 63828 382032
rect 39672 382016 39724 382022
rect 39672 381958 39724 381964
rect 24952 357944 25004 357950
rect 24952 357886 25004 357892
rect 24860 313404 24912 313410
rect 24860 313346 24912 313352
rect 24860 312792 24912 312798
rect 24860 312734 24912 312740
rect 24768 272128 24820 272134
rect 24768 272070 24820 272076
rect 24676 271992 24728 271998
rect 24676 271934 24728 271940
rect 24688 234705 24716 271934
rect 24674 234696 24730 234705
rect 24674 234631 24730 234640
rect 24780 199073 24808 272070
rect 24766 199064 24822 199073
rect 24766 198999 24822 199008
rect 24872 163441 24900 312734
rect 24858 163432 24914 163441
rect 24858 163367 24914 163376
rect 24964 128081 24992 357886
rect 147128 357808 147180 357814
rect 147128 357750 147180 357756
rect 122104 312928 122156 312934
rect 122104 312870 122156 312876
rect 98552 312860 98604 312866
rect 98552 312802 98604 312808
rect 98564 276758 98592 312802
rect 98000 276752 98052 276758
rect 98000 276694 98052 276700
rect 98552 276752 98604 276758
rect 98552 276694 98604 276700
rect 73896 276208 73948 276214
rect 73896 276150 73948 276156
rect 49976 276004 50028 276010
rect 49976 275946 50028 275952
rect 49988 273578 50016 275946
rect 73908 273578 73936 276150
rect 98012 273578 98040 276694
rect 122116 273578 122144 312870
rect 147140 276350 147168 357750
rect 268580 339998 268608 699858
rect 270500 627156 270552 627162
rect 270500 627098 270552 627104
rect 270408 586152 270460 586158
rect 270408 586094 270460 586100
rect 268842 512000 268898 512009
rect 268842 511935 268898 511944
rect 268856 510950 268884 511935
rect 268844 510944 268896 510950
rect 268844 510886 268896 510892
rect 270040 472592 270092 472598
rect 270040 472534 270092 472540
rect 269302 440736 269358 440745
rect 269302 440671 269358 440680
rect 269316 440162 269344 440671
rect 269304 440156 269356 440162
rect 269304 440098 269356 440104
rect 269302 405376 269358 405385
rect 269302 405311 269358 405320
rect 269316 404870 269344 405311
rect 269304 404864 269356 404870
rect 269304 404806 269356 404812
rect 269856 353252 269908 353258
rect 269856 353194 269908 353200
rect 269868 350334 269896 353194
rect 269856 350328 269908 350334
rect 269856 350270 269908 350276
rect 270052 348809 270080 472534
rect 270132 382356 270184 382362
rect 270132 382298 270184 382304
rect 270144 382090 270172 382298
rect 270132 382084 270184 382090
rect 270132 382026 270184 382032
rect 270144 353258 270172 382026
rect 270316 354068 270368 354074
rect 270316 354010 270368 354016
rect 270222 353832 270278 353841
rect 270222 353767 270278 353776
rect 270132 353252 270184 353258
rect 270132 353194 270184 353200
rect 270038 348800 270094 348809
rect 270038 348735 270094 348744
rect 269948 340060 270000 340066
rect 269948 340002 270000 340008
rect 268568 339992 268620 339998
rect 268568 339934 268620 339940
rect 269672 339992 269724 339998
rect 269960 339969 269988 340002
rect 269672 339934 269724 339940
rect 269946 339960 270002 339969
rect 269684 339697 269712 339934
rect 269946 339895 270002 339904
rect 270130 339824 270186 339833
rect 270130 339759 270186 339768
rect 269670 339688 269726 339697
rect 269670 339623 269726 339632
rect 270144 335617 270172 339759
rect 269854 335608 269910 335617
rect 269854 335543 269910 335552
rect 270130 335608 270186 335617
rect 270130 335543 270186 335552
rect 269394 329896 269450 329905
rect 269394 329831 269450 329840
rect 269408 329798 269436 329831
rect 268568 329792 268620 329798
rect 268568 329734 268620 329740
rect 269396 329792 269448 329798
rect 269396 329734 269448 329740
rect 146208 276344 146260 276350
rect 146208 276286 146260 276292
rect 147128 276344 147180 276350
rect 147128 276286 147180 276292
rect 146220 273578 146248 276286
rect 237012 276208 237064 276214
rect 237010 276176 237012 276185
rect 247224 276208 247276 276214
rect 237064 276176 237066 276185
rect 170128 276140 170180 276146
rect 170128 276082 170180 276088
rect 194232 276140 194284 276146
rect 237010 276111 237066 276120
rect 247222 276176 247224 276185
rect 247276 276176 247278 276185
rect 247222 276111 247278 276120
rect 194232 276082 194284 276088
rect 170140 273578 170168 276082
rect 194244 273578 194272 276082
rect 218336 276072 218388 276078
rect 218336 276014 218388 276020
rect 218348 273578 218376 276014
rect 242440 275392 242492 275398
rect 242440 275334 242492 275340
rect 242452 273578 242480 275334
rect 266360 275324 266412 275330
rect 266360 275266 266412 275272
rect 266372 273578 266400 275266
rect 49680 273550 50016 273578
rect 73600 273550 73936 273578
rect 97704 273550 98040 273578
rect 121808 273550 122144 273578
rect 145912 273550 146248 273578
rect 169832 273550 170168 273578
rect 193936 273550 194272 273578
rect 218040 273550 218376 273578
rect 242144 273550 242480 273578
rect 266064 273550 266400 273578
rect 27252 272400 27304 272406
rect 27252 272342 27304 272348
rect 27264 270881 27292 272342
rect 27250 270872 27306 270881
rect 27250 270807 27306 270816
rect 268384 238468 268436 238474
rect 268384 238410 268436 238416
rect 268396 237425 268424 238410
rect 268382 237416 268438 237425
rect 268382 237351 268438 237360
rect 268384 202836 268436 202842
rect 268384 202778 268436 202784
rect 268396 201793 268424 202778
rect 268382 201784 268438 201793
rect 268382 201719 268438 201728
rect 268580 166161 268608 329734
rect 269868 322402 269896 335543
rect 269868 322374 270080 322402
rect 270052 312186 270080 322374
rect 270040 312180 270092 312186
rect 270040 312122 270092 312128
rect 270040 312044 270092 312050
rect 270040 311986 270092 311992
rect 270052 309126 270080 311986
rect 270040 309120 270092 309126
rect 270040 309062 270092 309068
rect 269856 297424 269908 297430
rect 269856 297366 269908 297372
rect 269868 293350 269896 297366
rect 269856 293344 269908 293350
rect 269856 293286 269908 293292
rect 269948 287088 270000 287094
rect 269948 287030 270000 287036
rect 269960 260522 269988 287030
rect 270236 276078 270264 353767
rect 270328 324465 270356 354010
rect 270420 345273 270448 586094
rect 270406 345264 270462 345273
rect 270406 345199 270462 345208
rect 270314 324456 270370 324465
rect 270314 324391 270370 324400
rect 270420 276146 270448 345199
rect 270512 320793 270540 627098
rect 270592 586152 270644 586158
rect 270592 586094 270644 586100
rect 270604 586022 270632 586094
rect 270592 586016 270644 586022
rect 270592 585958 270644 585964
rect 270604 353841 270632 585958
rect 270590 353832 270646 353841
rect 270590 353767 270646 353776
rect 270590 350840 270646 350849
rect 270590 350775 270646 350784
rect 270498 320784 270554 320793
rect 270498 320719 270554 320728
rect 270408 276140 270460 276146
rect 270408 276082 270460 276088
rect 270224 276072 270276 276078
rect 270224 276014 270276 276020
rect 269960 260494 270080 260522
rect 270052 250322 270080 260494
rect 270052 250294 270264 250322
rect 270144 237046 270172 237077
rect 270236 237046 270264 250294
rect 270132 237040 270184 237046
rect 270224 237040 270276 237046
rect 270222 237008 270224 237017
rect 270276 237008 270278 237017
rect 270184 236988 270222 236994
rect 270132 236982 270222 236988
rect 270144 236966 270222 236982
rect 270222 236943 270278 236952
rect 270406 237008 270462 237017
rect 270406 236943 270462 236952
rect 270420 226778 270448 236943
rect 270224 226772 270276 226778
rect 270224 226714 270276 226720
rect 270408 226772 270460 226778
rect 270408 226714 270460 226720
rect 270236 216442 270264 226714
rect 270132 216436 270184 216442
rect 270132 216378 270184 216384
rect 270224 216436 270276 216442
rect 270224 216378 270276 216384
rect 270144 216345 270172 216378
rect 270130 216336 270186 216345
rect 270130 216271 270186 216280
rect 270222 206136 270278 206145
rect 270222 206071 270278 206080
rect 270236 195906 270264 206071
rect 270224 195900 270276 195906
rect 270144 195838 270172 195869
rect 270224 195842 270276 195848
rect 270132 195832 270184 195838
rect 270222 195800 270278 195809
rect 270184 195780 270222 195786
rect 270132 195774 270222 195780
rect 270144 195758 270222 195774
rect 270222 195735 270278 195744
rect 270406 195800 270462 195809
rect 270406 195735 270462 195744
rect 270420 185570 270448 195735
rect 270224 185564 270276 185570
rect 270224 185506 270276 185512
rect 270408 185564 270460 185570
rect 270408 185506 270460 185512
rect 270236 185473 270264 185506
rect 269946 185464 270002 185473
rect 269946 185399 270002 185408
rect 270222 185464 270278 185473
rect 270222 185399 270278 185408
rect 269960 175234 269988 185399
rect 269948 175228 270000 175234
rect 269948 175170 270000 175176
rect 270132 175228 270184 175234
rect 270132 175170 270184 175176
rect 270144 175114 270172 175170
rect 270222 175128 270278 175137
rect 270144 175086 270222 175114
rect 270222 175063 270278 175072
rect 270406 175128 270462 175137
rect 270406 175063 270462 175072
rect 268566 166152 268622 166161
rect 268566 166087 268622 166096
rect 270420 164898 270448 175063
rect 270224 164892 270276 164898
rect 270224 164834 270276 164840
rect 270408 164892 270460 164898
rect 270408 164834 270460 164840
rect 270236 164801 270264 164834
rect 270222 164792 270278 164801
rect 270222 164727 270278 164736
rect 270406 164792 270462 164801
rect 270406 164727 270462 164736
rect 270420 157486 270448 164727
rect 270132 157480 270184 157486
rect 270132 157422 270184 157428
rect 270408 157480 270460 157486
rect 270408 157422 270460 157428
rect 270144 152930 270172 157422
rect 270132 152924 270184 152930
rect 270132 152866 270184 152872
rect 270224 144288 270276 144294
rect 270144 144236 270224 144242
rect 270144 144230 270276 144236
rect 270144 144214 270264 144230
rect 270144 134065 270172 144214
rect 270130 134056 270186 134065
rect 270130 133991 270186 134000
rect 270130 132560 270186 132569
rect 270130 132495 270186 132504
rect 270144 131034 270172 132495
rect 270132 131028 270184 131034
rect 270132 130970 270184 130976
rect 267922 130520 267978 130529
rect 267922 130455 267978 130464
rect 267936 130286 267964 130455
rect 267924 130280 267976 130286
rect 267924 130222 267976 130228
rect 24950 128072 25006 128081
rect 24950 128007 25006 128016
rect 270224 120760 270276 120766
rect 270224 120702 270276 120708
rect 270236 116346 270264 120702
rect 270224 116340 270276 116346
rect 270224 116282 270276 116288
rect 270316 116204 270368 116210
rect 270316 116146 270368 116152
rect 270328 101658 270356 116146
rect 270224 101652 270276 101658
rect 270224 101594 270276 101600
rect 270316 101652 270368 101658
rect 270316 101594 270368 101600
rect 270236 101538 270264 101594
rect 270144 101510 270264 101538
rect 267922 95160 267978 95169
rect 267922 95095 267978 95104
rect 267936 94926 267964 95095
rect 267924 94920 267976 94926
rect 267924 94862 267976 94868
rect 24950 92440 25006 92449
rect 24950 92375 25006 92384
rect 24964 76022 24992 92375
rect 270144 91322 270172 101510
rect 270040 91316 270092 91322
rect 270040 91258 270092 91264
rect 270132 91316 270184 91322
rect 270132 91258 270184 91264
rect 270052 85490 270080 91258
rect 269960 85462 270080 85490
rect 269960 82414 269988 85462
rect 269672 82408 269724 82414
rect 269672 82350 269724 82356
rect 269948 82408 270000 82414
rect 269948 82350 270000 82356
rect 24952 76016 25004 76022
rect 24952 75958 25004 75964
rect 39376 73630 39712 73658
rect 63480 73630 63816 73658
rect 87400 73630 87736 73658
rect 111504 73630 111840 73658
rect 135608 73630 135944 73658
rect 159712 73630 160048 73658
rect 183816 73630 183968 73658
rect 207736 73630 208072 73658
rect 231840 73630 232176 73658
rect 255944 73630 256096 73658
rect 39684 72078 39712 73630
rect 39672 72072 39724 72078
rect 39672 72014 39724 72020
rect 63788 71602 63816 73630
rect 87708 72010 87736 73630
rect 87696 72004 87748 72010
rect 87696 71946 87748 71952
rect 111812 71806 111840 73630
rect 135916 71874 135944 73630
rect 160020 71942 160048 73630
rect 160008 71936 160060 71942
rect 160008 71878 160060 71884
rect 135904 71868 135956 71874
rect 135904 71810 135956 71816
rect 111800 71800 111852 71806
rect 111800 71742 111852 71748
rect 183940 71738 183968 73630
rect 183928 71732 183980 71738
rect 183928 71674 183980 71680
rect 208044 71670 208072 73630
rect 208032 71664 208084 71670
rect 208032 71606 208084 71612
rect 63776 71596 63828 71602
rect 63776 71538 63828 71544
rect 232148 71534 232176 73630
rect 256068 72146 256096 73630
rect 269684 72185 269712 82350
rect 269670 72176 269726 72185
rect 256056 72140 256108 72146
rect 269670 72111 269726 72120
rect 269854 72176 269910 72185
rect 269854 72111 269910 72120
rect 256056 72082 256108 72088
rect 269868 72026 269896 72111
rect 269776 71998 269896 72026
rect 269776 71602 269804 71998
rect 269764 71596 269816 71602
rect 269764 71538 269816 71544
rect 232136 71528 232188 71534
rect 232136 71470 232188 71476
rect 270604 3670 270632 350775
rect 270696 333713 270724 699926
rect 270776 699916 270828 699922
rect 270776 699858 270828 699864
rect 270682 333704 270738 333713
rect 270682 333639 270738 333648
rect 270788 317801 270816 699858
rect 271880 575544 271932 575550
rect 271880 575486 271932 575492
rect 271892 571266 271920 575486
rect 271880 571260 271932 571266
rect 271880 571202 271932 571208
rect 272340 382560 272392 382566
rect 272340 382502 272392 382508
rect 272352 381993 272380 382502
rect 272338 381984 272394 381993
rect 272338 381919 272394 381928
rect 272996 343058 273024 700062
rect 273076 700052 273128 700058
rect 273076 699994 273128 700000
rect 272984 343052 273036 343058
rect 272984 342994 273036 343000
rect 273088 342530 273116 699994
rect 273536 359236 273588 359242
rect 273536 359178 273588 359184
rect 273168 357876 273220 357882
rect 273168 357818 273220 357824
rect 272996 342502 273116 342530
rect 272996 342446 273024 342502
rect 272616 342440 272668 342446
rect 272614 342408 272616 342417
rect 272984 342440 273036 342446
rect 272668 342408 272670 342417
rect 272984 342382 273036 342388
rect 272614 342343 272670 342352
rect 272892 340060 272944 340066
rect 272892 340002 272944 340008
rect 272904 332738 272932 340002
rect 272904 332710 273116 332738
rect 272614 327584 272670 327593
rect 273088 327570 273116 332710
rect 272670 327542 273116 327570
rect 272614 327519 272670 327528
rect 270774 317792 270830 317801
rect 270774 317727 270830 317736
rect 273180 71942 273208 357818
rect 273548 71942 273576 359178
rect 273824 355586 273852 700606
rect 283852 700126 283880 703520
rect 332520 700670 332548 703520
rect 332508 700664 332560 700670
rect 332508 700606 332560 700612
rect 283840 700120 283892 700126
rect 283840 700062 283892 700068
rect 364996 700058 365024 703520
rect 397472 700670 397500 703520
rect 397460 700664 397512 700670
rect 397460 700606 397512 700612
rect 364984 700052 365036 700058
rect 364984 699994 365036 700000
rect 429856 699990 429884 703520
rect 462332 700670 462360 703520
rect 462320 700664 462372 700670
rect 462320 700606 462372 700612
rect 429844 699984 429896 699990
rect 494808 699961 494836 703520
rect 527192 700670 527220 703520
rect 527180 700664 527232 700670
rect 527180 700606 527232 700612
rect 527192 699990 527220 700606
rect 527180 699984 527232 699990
rect 429844 699926 429896 699932
rect 494794 699952 494850 699961
rect 527180 699926 527232 699932
rect 559668 699922 559696 703520
rect 579896 699984 579948 699990
rect 579896 699926 579948 699932
rect 494794 699887 494850 699896
rect 559656 699916 559708 699922
rect 559656 699858 559708 699864
rect 579908 698057 579936 699926
rect 579894 698048 579950 698057
rect 579894 697983 579950 697992
rect 579158 674656 579214 674665
rect 579158 674591 579214 674600
rect 578790 627736 578846 627745
rect 578790 627671 578846 627680
rect 578804 627162 578832 627671
rect 578792 627156 578844 627162
rect 578792 627098 578844 627104
rect 307574 586528 307630 586537
rect 307574 586463 307576 586472
rect 307628 586463 307630 586472
rect 341522 586528 341578 586537
rect 341522 586463 341578 586472
rect 485780 586492 485832 586498
rect 307576 586434 307628 586440
rect 289452 586424 289504 586430
rect 289450 586392 289452 586401
rect 289504 586392 289506 586401
rect 289450 586327 289506 586336
rect 293592 586356 293644 586362
rect 289464 586129 289492 586327
rect 293592 586298 293644 586304
rect 289450 586120 289506 586129
rect 284760 586084 284812 586090
rect 293604 586090 293632 586298
rect 298652 586288 298704 586294
rect 298652 586230 298704 586236
rect 298664 586129 298692 586230
rect 298650 586120 298706 586129
rect 289450 586055 289506 586064
rect 293592 586084 293644 586090
rect 284760 586026 284812 586032
rect 298650 586055 298706 586064
rect 293592 586026 293644 586032
rect 276664 582344 276716 582350
rect 276664 582286 276716 582292
rect 276676 580718 276704 582286
rect 276664 580712 276716 580718
rect 276664 580654 276716 580660
rect 276572 571124 276624 571130
rect 276572 571066 276624 571072
rect 276584 566710 276612 571066
rect 276572 566704 276624 566710
rect 276572 566646 276624 566652
rect 276388 510944 276440 510950
rect 276386 510912 276388 510921
rect 276440 510912 276442 510921
rect 276386 510847 276442 510856
rect 273904 382696 273956 382702
rect 273904 382638 273956 382644
rect 273916 382265 273944 382638
rect 273902 382256 273958 382265
rect 273902 382191 273958 382200
rect 276676 356538 276704 580654
rect 279240 566704 279292 566710
rect 279240 566646 279292 566652
rect 279252 560114 279280 566646
rect 279240 560108 279292 560114
rect 279240 560050 279292 560056
rect 280344 560108 280396 560114
rect 280344 560050 280396 560056
rect 280356 538762 280384 560050
rect 280344 538756 280396 538762
rect 280344 538698 280396 538704
rect 282184 538756 282236 538762
rect 282184 538698 282236 538704
rect 282196 535090 282224 538698
rect 282184 535084 282236 535090
rect 282184 535026 282236 535032
rect 284116 516724 284168 516730
rect 284116 516666 284168 516672
rect 284128 515234 284156 516666
rect 283288 515228 283340 515234
rect 283288 515170 283340 515176
rect 284116 515228 284168 515234
rect 284116 515170 284168 515176
rect 283300 510921 283328 515170
rect 283286 510912 283342 510921
rect 283286 510847 283342 510856
rect 278228 382424 278280 382430
rect 278228 382366 278280 382372
rect 279608 382424 279660 382430
rect 279608 382366 279660 382372
rect 278240 373810 278268 382366
rect 279620 382090 279648 382366
rect 279700 382220 279752 382226
rect 279700 382162 279752 382168
rect 279608 382084 279660 382090
rect 279608 382026 279660 382032
rect 278240 373782 278360 373810
rect 278332 363610 278360 373782
rect 278332 363582 278544 363610
rect 278516 359242 278544 363582
rect 279712 359281 279740 382162
rect 279698 359272 279754 359281
rect 278504 359236 278556 359242
rect 279698 359207 279754 359216
rect 280618 359272 280674 359281
rect 280618 359207 280674 359216
rect 278504 359178 278556 359184
rect 276676 356510 276796 356538
rect 273824 355558 274036 355586
rect 274008 355450 274036 355558
rect 274008 355422 274390 355450
rect 276768 354929 276796 356510
rect 278516 355450 278544 359178
rect 278516 355422 278622 355450
rect 280632 355436 280660 359207
rect 284772 358494 284800 586026
rect 289176 585948 289228 585954
rect 289176 585890 289228 585896
rect 288532 535084 288584 535090
rect 288532 535026 288584 535032
rect 288544 534002 288572 535026
rect 288532 533996 288584 534002
rect 288532 533938 288584 533944
rect 287060 523252 287112 523258
rect 287060 523194 287112 523200
rect 287072 519738 287100 523194
rect 286980 519710 287100 519738
rect 286980 516730 287008 519710
rect 286968 516724 287020 516730
rect 286968 516666 287020 516672
rect 286232 440156 286284 440162
rect 286232 440098 286284 440104
rect 286244 386306 286272 440098
rect 286232 386300 286284 386306
rect 286232 386242 286284 386248
rect 286244 385762 286272 386242
rect 286232 385756 286284 385762
rect 286232 385698 286284 385704
rect 286692 385756 286744 385762
rect 286692 385698 286744 385704
rect 284760 358488 284812 358494
rect 284760 358430 284812 358436
rect 282644 358420 282696 358426
rect 282644 358362 282696 358368
rect 282656 355436 282684 358362
rect 284668 357808 284720 357814
rect 284668 357750 284720 357756
rect 284680 355436 284708 357750
rect 276754 354920 276810 354929
rect 276598 354878 276754 354906
rect 286704 354906 286732 385698
rect 289188 354929 289216 585890
rect 290004 533996 290056 534002
rect 290004 533938 290056 533944
rect 289268 528488 289320 528494
rect 289268 528430 289320 528436
rect 289280 523258 289308 528430
rect 290016 526998 290044 533938
rect 291384 533724 291436 533730
rect 291384 533666 291436 533672
rect 291396 528494 291424 533666
rect 291384 528488 291436 528494
rect 291384 528430 291436 528436
rect 290004 526992 290056 526998
rect 290004 526934 290056 526940
rect 292764 526992 292816 526998
rect 292764 526934 292816 526940
rect 292776 524074 292804 526934
rect 292764 524068 292816 524074
rect 292764 524010 292816 524016
rect 289268 523252 289320 523258
rect 289268 523194 289320 523200
rect 293604 354929 293632 586026
rect 300216 586016 300268 586022
rect 300216 585958 300268 585964
rect 299572 554396 299624 554402
rect 299572 554338 299624 554344
rect 299584 552090 299612 554338
rect 297364 552084 297416 552090
rect 297364 552026 297416 552032
rect 299572 552084 299624 552090
rect 299572 552026 299624 552032
rect 297376 543794 297404 552026
rect 295892 543788 295944 543794
rect 295892 543730 295944 543736
rect 297364 543788 297416 543794
rect 297364 543730 297416 543736
rect 295904 538082 295932 543730
rect 294420 538076 294472 538082
rect 294420 538018 294472 538024
rect 295892 538076 295944 538082
rect 295892 538018 295944 538024
rect 294432 533730 294460 538018
rect 294420 533724 294472 533730
rect 294420 533666 294472 533672
rect 295524 524000 295576 524006
rect 295524 523942 295576 523948
rect 295536 521082 295564 523942
rect 295524 521076 295576 521082
rect 295524 521018 295576 521024
rect 298468 521076 298520 521082
rect 298468 521018 298520 521024
rect 298480 516730 298508 521018
rect 298468 516724 298520 516730
rect 298468 516666 298520 516672
rect 297272 382628 297324 382634
rect 297272 382570 297324 382576
rect 297284 382129 297312 382570
rect 297270 382120 297326 382129
rect 297270 382055 297326 382064
rect 300228 358902 300256 585958
rect 341536 583930 341564 586463
rect 485780 586434 485832 586440
rect 365442 586392 365498 586401
rect 365442 586327 365498 586336
rect 365456 583930 365484 586327
rect 413650 586256 413706 586265
rect 413650 586191 413706 586200
rect 413664 583930 413692 586191
rect 461674 586120 461730 586129
rect 461674 586055 461730 586064
rect 437756 586016 437808 586022
rect 437756 585958 437808 585964
rect 437768 583930 437796 585958
rect 461688 583930 461716 586055
rect 485792 583930 485820 586434
rect 509884 586152 509936 586158
rect 509884 586094 509936 586100
rect 509896 583930 509924 586094
rect 533988 586084 534040 586090
rect 533988 586026 534040 586032
rect 534000 583930 534028 586026
rect 557908 585948 557960 585954
rect 557908 585890 557960 585896
rect 557920 583930 557948 585890
rect 341536 583902 341826 583930
rect 365456 583902 365746 583930
rect 413664 583902 413954 583930
rect 437768 583902 438058 583930
rect 461688 583902 461978 583930
rect 485792 583902 486082 583930
rect 509896 583902 510186 583930
rect 534000 583902 534290 583930
rect 557920 583902 558210 583930
rect 314384 582480 314436 582486
rect 314384 582422 314436 582428
rect 313464 582276 313516 582282
rect 313464 582218 313516 582224
rect 309140 574048 309192 574054
rect 309140 573990 309192 573996
rect 309152 571878 309180 573990
rect 305368 571872 305420 571878
rect 305368 571814 305420 571820
rect 309140 571872 309192 571878
rect 309140 571814 309192 571820
rect 305380 557938 305408 571814
rect 305368 557932 305420 557938
rect 305368 557874 305420 557880
rect 301688 557864 301740 557870
rect 301688 557806 301740 557812
rect 301700 554402 301728 557806
rect 301688 554396 301740 554402
rect 301688 554338 301740 554344
rect 313476 549030 313504 582218
rect 314396 565282 314424 582422
rect 319444 582344 319496 582350
rect 319444 582286 319496 582292
rect 558736 582344 558788 582350
rect 558736 582286 558788 582292
rect 315396 580712 315448 580718
rect 315394 580680 315396 580689
rect 315448 580680 315450 580689
rect 315394 580615 315450 580624
rect 319456 578542 319484 582286
rect 558552 580032 558604 580038
rect 558552 579974 558604 579980
rect 317972 578536 318024 578542
rect 317972 578478 318024 578484
rect 319444 578536 319496 578542
rect 319444 578478 319496 578484
rect 317984 574122 318012 578478
rect 317972 574116 318024 574122
rect 317972 574058 318024 574064
rect 314108 565276 314160 565282
rect 314108 565218 314160 565224
rect 314384 565276 314436 565282
rect 314384 565218 314436 565224
rect 314120 565185 314148 565218
rect 314106 565176 314162 565185
rect 314106 565111 314162 565120
rect 314198 559328 314254 559337
rect 314198 559263 314254 559272
rect 314212 549114 314240 559263
rect 314120 549086 314240 549114
rect 313464 549024 313516 549030
rect 313464 548966 313516 548972
rect 314120 548978 314148 549086
rect 313476 547670 313504 548966
rect 314120 548950 314240 548978
rect 313464 547664 313516 547670
rect 313464 547606 313516 547612
rect 313924 547664 313976 547670
rect 313924 547606 313976 547612
rect 301780 516724 301832 516730
rect 301780 516666 301832 516672
rect 301792 513806 301820 516666
rect 301780 513800 301832 513806
rect 301780 513742 301832 513748
rect 306104 513732 306156 513738
rect 306104 513674 306156 513680
rect 306116 510898 306144 513674
rect 306116 510870 306236 510898
rect 306208 509726 306236 510870
rect 306196 509720 306248 509726
rect 306196 509662 306248 509668
rect 307576 509720 307628 509726
rect 307576 509662 307628 509668
rect 303896 404864 303948 404870
rect 303896 404806 303948 404812
rect 303908 385665 303936 404806
rect 303894 385656 303950 385665
rect 303894 385591 303950 385600
rect 300952 382424 301004 382430
rect 300952 382366 301004 382372
rect 300964 382022 300992 382366
rect 300952 382016 301004 382022
rect 300952 381958 301004 381964
rect 299020 358896 299072 358902
rect 299020 358838 299072 358844
rect 300216 358896 300268 358902
rect 300216 358838 300268 358844
rect 294972 358488 295024 358494
rect 294972 358430 295024 358436
rect 294984 355436 295012 358430
rect 296996 357876 297048 357882
rect 296996 357818 297048 357824
rect 297008 355436 297036 357818
rect 299032 355436 299060 358838
rect 300964 354929 300992 381958
rect 305276 358556 305328 358562
rect 305276 358498 305328 358504
rect 303252 358488 303304 358494
rect 303252 358430 303304 358436
rect 303264 355436 303292 358430
rect 305288 355436 305316 358498
rect 286966 354920 287022 354929
rect 286704 354892 286966 354906
rect 286718 354878 286966 354892
rect 276754 354855 276810 354864
rect 289174 354920 289230 354929
rect 288926 354878 289174 354906
rect 286966 354855 287022 354864
rect 291198 354920 291254 354929
rect 290950 354878 291198 354906
rect 289174 354855 289230 354864
rect 293222 354920 293278 354929
rect 292974 354878 293222 354906
rect 291198 354855 291254 354864
rect 293222 354855 293278 354864
rect 293590 354920 293646 354929
rect 293590 354855 293646 354864
rect 300950 354920 301006 354929
rect 306930 354920 306986 354929
rect 301006 354878 301254 354906
rect 300950 354855 301006 354864
rect 307588 354906 307616 509662
rect 313740 386368 313792 386374
rect 313740 386310 313792 386316
rect 313648 382288 313700 382294
rect 313648 382230 313700 382236
rect 311348 357944 311400 357950
rect 311348 357886 311400 357892
rect 311360 355436 311388 357886
rect 306986 354878 307616 354906
rect 309350 354890 309640 354906
rect 309350 354884 309652 354890
rect 309350 354878 309600 354884
rect 306930 354855 306986 354864
rect 309600 354826 309652 354832
rect 312728 354884 312780 354890
rect 312728 354826 312780 354832
rect 311532 354136 311584 354142
rect 311532 354078 311584 354084
rect 311544 352073 311572 354078
rect 311530 352064 311586 352073
rect 311530 351999 311586 352008
rect 296534 316296 296590 316305
rect 296286 316254 296534 316282
rect 298558 316296 298614 316305
rect 296534 316231 296590 316240
rect 298020 316254 298558 316282
rect 294262 315846 294460 315874
rect 281184 315710 281934 315738
rect 275926 315616 275982 315625
rect 275678 315588 275926 315602
rect 273640 313410 273668 315588
rect 275664 315574 275926 315588
rect 273628 313404 273680 313410
rect 273628 313346 273680 313352
rect 275664 312769 275692 315574
rect 275926 315551 275982 315560
rect 277688 313449 277716 315588
rect 279712 315574 279910 315602
rect 277674 313440 277730 313449
rect 277674 313375 277730 313384
rect 279712 313177 279740 315574
rect 281184 313313 281212 315710
rect 281170 313304 281226 313313
rect 283944 313290 283972 315588
rect 285968 313478 285996 315588
rect 285956 313472 286008 313478
rect 285956 313414 286008 313420
rect 287992 313410 288020 315588
rect 287980 313404 288032 313410
rect 287980 313346 288032 313352
rect 284022 313304 284078 313313
rect 283944 313262 284022 313290
rect 281170 313239 281226 313248
rect 284022 313239 284078 313248
rect 279698 313168 279754 313177
rect 279698 313103 279754 313112
rect 275650 312760 275706 312769
rect 275650 312695 275706 312704
rect 276570 312760 276626 312769
rect 276570 312695 276626 312704
rect 276584 272066 276612 312695
rect 276662 273728 276718 273737
rect 276662 273663 276718 273672
rect 276676 272406 276704 273663
rect 276664 272400 276716 272406
rect 276664 272342 276716 272348
rect 276572 272060 276624 272066
rect 276572 272002 276624 272008
rect 276584 271794 276612 272002
rect 275928 271788 275980 271794
rect 275928 271730 275980 271736
rect 276572 271788 276624 271794
rect 276572 271730 276624 271736
rect 275940 202842 275968 271730
rect 276676 270842 276704 272342
rect 276664 270836 276716 270842
rect 276664 270778 276716 270784
rect 275928 202836 275980 202842
rect 275928 202778 275980 202784
rect 279712 72146 279740 313103
rect 279700 72140 279752 72146
rect 279700 72082 279752 72088
rect 276662 72040 276718 72049
rect 281184 72010 281212 313239
rect 284036 276350 284064 313239
rect 290016 312934 290044 315588
rect 292224 313478 292252 315588
rect 292212 313472 292264 313478
rect 292212 313414 292264 313420
rect 290004 312928 290056 312934
rect 290004 312870 290056 312876
rect 294432 312338 294460 315846
rect 294340 312310 294460 312338
rect 289818 276720 289874 276729
rect 289818 276655 289874 276664
rect 293590 276720 293646 276729
rect 293590 276655 293646 276664
rect 284024 276344 284076 276350
rect 284024 276286 284076 276292
rect 284036 276214 284064 276286
rect 284024 276208 284076 276214
rect 284024 276150 284076 276156
rect 289832 275330 289860 276655
rect 293604 275398 293632 276655
rect 294340 276350 294368 312310
rect 294328 276344 294380 276350
rect 294328 276286 294380 276292
rect 293592 275392 293644 275398
rect 293592 275334 293644 275340
rect 289820 275324 289872 275330
rect 289820 275266 289872 275272
rect 286230 133920 286286 133929
rect 286230 133855 286286 133864
rect 286244 130286 286272 133855
rect 286232 130280 286284 130286
rect 286232 130222 286284 130228
rect 286244 114850 286272 130222
rect 286232 114844 286284 114850
rect 286232 114786 286284 114792
rect 289544 114776 289596 114782
rect 289544 114718 289596 114724
rect 289556 111858 289584 114718
rect 289544 111852 289596 111858
rect 289544 111794 289596 111800
rect 292856 111852 292908 111858
rect 292856 111794 292908 111800
rect 292868 109954 292896 111794
rect 292856 109948 292908 109954
rect 292856 109890 292908 109896
rect 294420 109948 294472 109954
rect 294420 109890 294472 109896
rect 294432 108934 294460 109890
rect 294420 108928 294472 108934
rect 294420 108870 294472 108876
rect 296548 72010 296576 316231
rect 298020 276214 298048 316254
rect 310886 316296 310942 316305
rect 310638 316254 310886 316282
rect 298558 316231 298614 316240
rect 310886 316231 310942 316240
rect 306746 315616 306802 315625
rect 300320 312866 300348 315588
rect 300308 312860 300360 312866
rect 300308 312802 300360 312808
rect 302528 312798 302556 315588
rect 304552 315489 304580 315588
rect 306590 315574 306746 315602
rect 306802 315574 306880 315602
rect 306746 315551 306802 315560
rect 306760 315491 306788 315551
rect 304538 315480 304594 315489
rect 304538 315415 304594 315424
rect 302516 312792 302568 312798
rect 304552 312769 304580 315415
rect 302516 312734 302568 312740
rect 303250 312760 303306 312769
rect 303250 312695 303306 312704
rect 304538 312760 304594 312769
rect 304538 312695 304594 312704
rect 298008 276208 298060 276214
rect 298008 276150 298060 276156
rect 297272 108928 297324 108934
rect 297272 108870 297324 108876
rect 297284 103034 297312 108870
rect 297284 103006 297404 103034
rect 297376 97646 297404 103006
rect 297364 97640 297416 97646
rect 297364 97582 297416 97588
rect 298836 97640 298888 97646
rect 298836 97582 298888 97588
rect 298848 89826 298876 97582
rect 303264 94926 303292 312695
rect 306852 276010 306880 315574
rect 308600 313546 308628 315588
rect 308588 313540 308640 313546
rect 308588 313482 308640 313488
rect 306840 276004 306892 276010
rect 306840 275946 306892 275952
rect 306838 272232 306894 272241
rect 306838 272167 306894 272176
rect 306852 272134 306880 272167
rect 306840 272128 306892 272134
rect 306840 272070 306892 272076
rect 306852 200190 306880 272070
rect 306840 200184 306892 200190
rect 306840 200126 306892 200132
rect 312740 164830 312768 354826
rect 313556 354000 313608 354006
rect 313556 353942 313608 353948
rect 313568 339969 313596 353942
rect 313554 339960 313610 339969
rect 313554 339895 313610 339904
rect 313554 330984 313610 330993
rect 313554 330919 313610 330928
rect 312728 164824 312780 164830
rect 312728 164766 312780 164772
rect 303252 94920 303304 94926
rect 303252 94862 303304 94868
rect 303896 94920 303948 94926
rect 303896 94862 303948 94868
rect 298836 89820 298888 89826
rect 298836 89762 298888 89768
rect 301780 89752 301832 89758
rect 301780 89694 301832 89700
rect 301792 86970 301820 89694
rect 301780 86964 301832 86970
rect 301780 86906 301832 86912
rect 303908 75954 303936 94862
rect 308956 86828 309008 86834
rect 308956 86770 309008 86776
rect 308968 84250 308996 86770
rect 308956 84244 309008 84250
rect 308956 84186 309008 84192
rect 312084 84244 312136 84250
rect 312084 84186 312136 84192
rect 312096 80986 312124 84186
rect 312084 80980 312136 80986
rect 312084 80922 312136 80928
rect 303896 75948 303948 75954
rect 303896 75890 303948 75896
rect 300952 72072 301004 72078
rect 300950 72040 300952 72049
rect 301004 72040 301006 72049
rect 276662 71975 276718 71984
rect 281172 72004 281224 72010
rect 273168 71936 273220 71942
rect 273168 71878 273220 71884
rect 273260 71936 273312 71942
rect 273260 71878 273312 71884
rect 273536 71936 273588 71942
rect 273536 71878 273588 71884
rect 273272 71670 273300 71878
rect 276676 71806 276704 71975
rect 281172 71946 281224 71952
rect 296076 72004 296128 72010
rect 296076 71946 296128 71952
rect 296536 72004 296588 72010
rect 300950 71975 301006 71984
rect 296536 71946 296588 71952
rect 276664 71800 276716 71806
rect 276664 71742 276716 71748
rect 281184 71670 281212 71946
rect 273260 71664 273312 71670
rect 273260 71606 273312 71612
rect 281172 71664 281224 71670
rect 281172 71606 281224 71612
rect 296088 71534 296116 71946
rect 300964 71534 300992 71975
rect 313568 71874 313596 330919
rect 313660 327593 313688 382230
rect 313752 345817 313780 386310
rect 313832 382152 313884 382158
rect 313832 382094 313884 382100
rect 313738 345808 313794 345817
rect 313738 345743 313794 345752
rect 313738 336560 313794 336569
rect 313738 336495 313794 336504
rect 313646 327584 313702 327593
rect 313646 327519 313702 327528
rect 313660 72078 313688 327519
rect 313752 271998 313780 336495
rect 313844 330993 313872 382094
rect 313936 348809 313964 547606
rect 314212 544882 314240 548950
rect 315854 544912 315910 544921
rect 314200 544876 314252 544882
rect 315854 544847 315856 544856
rect 314200 544818 314252 544824
rect 315908 544847 315910 544856
rect 315856 544818 315908 544824
rect 314212 538778 314240 544818
rect 314212 538750 314516 538778
rect 314488 522617 314516 538750
rect 314106 522608 314162 522617
rect 314106 522543 314162 522552
rect 314474 522608 314530 522617
rect 314474 522543 314530 522552
rect 314120 518242 314148 522543
rect 314120 518214 314332 518242
rect 314304 512310 314332 518214
rect 314292 512304 314344 512310
rect 314292 512246 314344 512252
rect 314568 512304 314620 512310
rect 314568 512246 314620 512252
rect 314580 504937 314608 512246
rect 315488 509720 315540 509726
rect 315488 509662 315540 509668
rect 315500 509561 315528 509662
rect 315486 509552 315542 509561
rect 315486 509487 315542 509496
rect 314382 504928 314438 504937
rect 314304 504898 314382 504914
rect 314292 504892 314382 504898
rect 314344 504886 314382 504892
rect 314382 504863 314438 504872
rect 314566 504928 314622 504937
rect 314566 504863 314622 504872
rect 314292 504834 314344 504840
rect 314384 494624 314436 494630
rect 314384 494566 314436 494572
rect 314396 487234 314424 494566
rect 314304 487206 314424 487234
rect 314304 484294 314332 487206
rect 314292 484288 314344 484294
rect 314292 484230 314344 484236
rect 314384 474020 314436 474026
rect 314384 473962 314436 473968
rect 314396 466562 314424 473962
rect 315486 473104 315542 473113
rect 315486 473039 315542 473048
rect 315500 472598 315528 473039
rect 315488 472592 315540 472598
rect 315488 472534 315540 472540
rect 314304 466534 314424 466562
rect 314304 463690 314332 466534
rect 314292 463684 314344 463690
rect 314292 463626 314344 463632
rect 314384 453416 314436 453422
rect 314384 453358 314436 453364
rect 314396 446026 314424 453358
rect 314304 445998 314424 446026
rect 314304 435810 314332 445998
rect 314292 435804 314344 435810
rect 314292 435746 314344 435752
rect 314384 435736 314436 435742
rect 314384 435678 314436 435684
rect 314396 432750 314424 435678
rect 314384 432744 314436 432750
rect 314384 432686 314436 432692
rect 314384 425400 314436 425406
rect 314384 425342 314436 425348
rect 314396 422498 314424 425342
rect 314396 422470 314516 422498
rect 314488 412214 314516 422470
rect 314292 412208 314344 412214
rect 314290 412176 314292 412185
rect 314476 412208 314528 412214
rect 314344 412176 314346 412185
rect 314476 412150 314528 412156
rect 314658 412176 314714 412185
rect 314290 412111 314346 412120
rect 314658 412111 314714 412120
rect 314672 401985 314700 412111
rect 316222 402112 316278 402121
rect 316222 402047 316278 402056
rect 314382 401976 314438 401985
rect 314200 401940 314252 401946
rect 314382 401911 314438 401920
rect 314658 401976 314714 401985
rect 316236 401946 316264 402047
rect 314658 401911 314714 401920
rect 316224 401940 316276 401946
rect 314200 401882 314252 401888
rect 314212 386374 314240 401882
rect 314396 394602 314424 401911
rect 316224 401882 316276 401888
rect 314384 394596 314436 394602
rect 314384 394538 314436 394544
rect 314384 394460 314436 394466
rect 314384 394402 314436 394408
rect 314200 386368 314252 386374
rect 314200 386310 314252 386316
rect 314396 384282 314424 394402
rect 314120 384254 314424 384282
rect 314120 384146 314148 384254
rect 314120 384118 314240 384146
rect 314212 373998 314240 384118
rect 331508 382430 331536 383996
rect 331496 382424 331548 382430
rect 331496 382366 331548 382372
rect 355612 382362 355640 383996
rect 355600 382356 355652 382362
rect 355600 382298 355652 382304
rect 314936 382288 314988 382294
rect 379532 382265 379560 383996
rect 314936 382230 314988 382236
rect 379518 382256 379574 382265
rect 314948 382022 314976 382230
rect 403636 382226 403664 383996
rect 379518 382191 379574 382200
rect 403624 382220 403676 382226
rect 403624 382162 403676 382168
rect 427740 382158 427768 383996
rect 427728 382152 427780 382158
rect 427728 382094 427780 382100
rect 475948 382022 475976 383996
rect 499868 382090 499896 383996
rect 523972 382129 524000 383996
rect 523958 382120 524014 382129
rect 499856 382084 499908 382090
rect 523958 382055 524014 382064
rect 499856 382026 499908 382032
rect 314936 382016 314988 382022
rect 314936 381958 314988 381964
rect 475936 382016 475988 382022
rect 548076 381993 548104 383996
rect 475936 381958 475988 381964
rect 548062 381984 548118 381993
rect 548062 381919 548118 381928
rect 314200 373992 314252 373998
rect 314200 373934 314252 373940
rect 314292 373924 314344 373930
rect 314292 373866 314344 373872
rect 314304 370977 314332 373866
rect 314106 370968 314162 370977
rect 314106 370903 314162 370912
rect 314290 370968 314346 370977
rect 314290 370903 314346 370912
rect 314120 360738 314148 370903
rect 314108 360732 314160 360738
rect 314108 360674 314160 360680
rect 314384 360732 314436 360738
rect 314384 360674 314436 360680
rect 314396 353394 314424 360674
rect 314384 353388 314436 353394
rect 314384 353330 314436 353336
rect 314292 353252 314344 353258
rect 314292 353194 314344 353200
rect 313922 348800 313978 348809
rect 313922 348735 313978 348744
rect 314198 345808 314254 345817
rect 314198 345743 314254 345752
rect 314108 343052 314160 343058
rect 314108 342994 314160 343000
rect 314120 336569 314148 342994
rect 314106 336560 314162 336569
rect 314106 336495 314162 336504
rect 313830 330984 313886 330993
rect 313830 330919 313886 330928
rect 313740 271992 313792 271998
rect 313740 271934 313792 271940
rect 313752 270910 313780 271934
rect 313740 270904 313792 270910
rect 313740 270846 313792 270852
rect 314212 92410 314240 345743
rect 314304 343058 314332 353194
rect 314382 348800 314438 348809
rect 314382 348735 314438 348744
rect 314292 343052 314344 343058
rect 314292 342994 314344 343000
rect 314396 272406 314424 348735
rect 558564 334150 558592 579974
rect 558644 532908 558696 532914
rect 558644 532850 558696 532856
rect 558656 358562 558684 532850
rect 558748 515166 558776 582286
rect 560852 582276 560904 582282
rect 560852 582218 560904 582224
rect 560864 547777 560892 582218
rect 578790 580816 578846 580825
rect 578790 580751 578846 580760
rect 578804 580038 578832 580751
rect 578792 580032 578844 580038
rect 578792 579974 578844 579980
rect 560850 547768 560906 547777
rect 560850 547703 560906 547712
rect 578790 533896 578846 533905
rect 578790 533831 578846 533840
rect 578804 532914 578832 533831
rect 578792 532908 578844 532914
rect 578792 532850 578844 532856
rect 558736 515160 558788 515166
rect 558736 515102 558788 515108
rect 559380 515160 559432 515166
rect 559380 515102 559432 515108
rect 559392 512145 559420 515102
rect 559378 512136 559434 512145
rect 559378 512071 559434 512080
rect 560850 440736 560906 440745
rect 560850 440671 560906 440680
rect 560864 437322 560892 440671
rect 560772 437294 560892 437322
rect 560772 432546 560800 437294
rect 558828 432540 558880 432546
rect 558828 432482 558880 432488
rect 560760 432540 560812 432546
rect 560760 432482 560812 432488
rect 558736 391604 558788 391610
rect 558736 391546 558788 391552
rect 558644 358556 558696 358562
rect 558644 358498 558696 358504
rect 314936 334144 314988 334150
rect 314936 334086 314988 334092
rect 558552 334144 558604 334150
rect 558552 334086 558604 334092
rect 314948 333849 314976 334086
rect 314934 333840 314990 333849
rect 314934 333775 314990 333784
rect 558748 313410 558776 391546
rect 558840 386306 558868 432482
rect 560850 405376 560906 405385
rect 560850 405311 560906 405320
rect 558828 386300 558880 386306
rect 558828 386242 558880 386248
rect 560864 385665 560892 405311
rect 578790 393000 578846 393009
rect 578790 392935 578846 392944
rect 578804 391610 578832 392935
rect 578792 391604 578844 391610
rect 578792 391546 578844 391552
rect 560850 385656 560906 385665
rect 560850 385591 560906 385600
rect 579172 313478 579200 674591
rect 579908 651137 579936 697983
rect 579894 651128 579950 651137
rect 579894 651063 579950 651072
rect 579908 604217 579936 651063
rect 579894 604208 579950 604217
rect 579894 604143 579950 604152
rect 579908 557297 579936 604143
rect 579894 557288 579950 557297
rect 579894 557223 579950 557232
rect 579908 510377 579936 557223
rect 579894 510368 579950 510377
rect 579894 510303 579950 510312
rect 579250 486840 579306 486849
rect 579250 486775 579306 486784
rect 579264 358494 579292 486775
rect 579908 463457 579936 510303
rect 579894 463448 579950 463457
rect 579894 463383 579950 463392
rect 579342 439920 579398 439929
rect 579342 439855 579398 439864
rect 579252 358488 579304 358494
rect 579252 358430 579304 358436
rect 579356 354074 579384 439855
rect 579908 419506 579936 463383
rect 579816 419478 579936 419506
rect 579816 416537 579844 419478
rect 579802 416528 579858 416537
rect 579802 416463 579858 416472
rect 579816 409306 579844 416463
rect 579448 409278 579844 409306
rect 579448 358426 579476 409278
rect 579436 358420 579488 358426
rect 579436 358362 579488 358368
rect 579344 354068 579396 354074
rect 579344 354010 579396 354016
rect 579160 313472 579212 313478
rect 579160 313414 579212 313420
rect 558736 313404 558788 313410
rect 558736 313346 558788 313352
rect 365720 276412 365772 276418
rect 365720 276354 365772 276360
rect 341800 276004 341852 276010
rect 341800 275946 341852 275952
rect 341812 273564 341840 275946
rect 365732 273564 365760 276354
rect 413928 276344 413980 276350
rect 413928 276286 413980 276292
rect 461952 276344 462004 276350
rect 461952 276286 462004 276292
rect 413940 273564 413968 276286
rect 438030 276040 438086 276049
rect 438030 275975 438086 275984
rect 438044 273564 438072 275975
rect 461964 273564 461992 276286
rect 486056 276140 486108 276146
rect 486056 276082 486108 276088
rect 486068 273564 486096 276082
rect 510160 276072 510212 276078
rect 510160 276014 510212 276020
rect 510172 273564 510200 276014
rect 534264 275392 534316 275398
rect 534264 275334 534316 275340
rect 534276 273564 534304 275334
rect 558184 275324 558236 275330
rect 558184 275266 558236 275272
rect 558196 273564 558224 275266
rect 314384 272400 314436 272406
rect 314384 272342 314436 272348
rect 560852 272400 560904 272406
rect 560852 272342 560904 272348
rect 314292 270904 314344 270910
rect 314292 270846 314344 270852
rect 314304 234705 314332 270846
rect 314396 238474 314424 272342
rect 558552 272060 558604 272066
rect 558552 272002 558604 272008
rect 315028 270836 315080 270842
rect 315028 270778 315080 270784
rect 315040 270337 315068 270778
rect 315026 270328 315082 270337
rect 315026 270263 315082 270272
rect 314384 238468 314436 238474
rect 314384 238410 314436 238416
rect 314290 234696 314346 234705
rect 314290 234631 314346 234640
rect 558564 206106 558592 272002
rect 560864 237425 560892 272342
rect 560850 237416 560906 237425
rect 560850 237351 560906 237360
rect 558552 206100 558604 206106
rect 558552 206042 558604 206048
rect 558920 206100 558972 206106
rect 558920 206042 558972 206048
rect 558932 201793 558960 206042
rect 558918 201784 558974 201793
rect 558918 201719 558974 201728
rect 315028 200184 315080 200190
rect 315028 200126 315080 200132
rect 315040 199073 315068 200126
rect 315026 199064 315082 199073
rect 315026 198999 315082 199008
rect 315028 164824 315080 164830
rect 315028 164766 315080 164772
rect 315040 163441 315068 164766
rect 315026 163432 315082 163441
rect 315026 163367 315082 163376
rect 559378 130520 559434 130529
rect 559378 130455 559434 130464
rect 559392 119270 559420 130455
rect 558552 119264 558604 119270
rect 558552 119206 558604 119212
rect 559380 119264 559432 119270
rect 559380 119206 559432 119212
rect 315026 92440 315082 92449
rect 314200 92404 314252 92410
rect 315026 92375 315028 92384
rect 314200 92346 314252 92352
rect 315080 92375 315082 92384
rect 315028 92346 315080 92352
rect 314212 76022 314240 92346
rect 316408 80980 316460 80986
rect 316408 80922 316460 80928
rect 316420 78010 316448 80922
rect 316420 77982 316540 78010
rect 316512 76022 316540 77982
rect 558564 76022 558592 119206
rect 560850 95160 560906 95169
rect 560850 95095 560906 95104
rect 314200 76016 314252 76022
rect 314200 75958 314252 75964
rect 316500 76016 316552 76022
rect 316500 75958 316552 75964
rect 558552 76016 558604 76022
rect 558552 75958 558604 75964
rect 560864 75954 560892 95095
rect 560852 75948 560904 75954
rect 560852 75890 560904 75896
rect 313648 72072 313700 72078
rect 313648 72014 313700 72020
rect 313556 71868 313608 71874
rect 313556 71810 313608 71816
rect 313660 71738 313688 72014
rect 313648 71732 313700 71738
rect 313648 71674 313700 71680
rect 331508 71534 331536 73644
rect 355612 71602 355640 73644
rect 379532 71670 379560 73644
rect 403636 71806 403664 73644
rect 427740 71874 427768 73644
rect 475948 72078 475976 73644
rect 475936 72072 475988 72078
rect 475936 72014 475988 72020
rect 499868 71942 499896 73644
rect 523972 72010 524000 73644
rect 548076 72146 548104 73644
rect 548064 72140 548116 72146
rect 548064 72082 548116 72088
rect 523960 72004 524012 72010
rect 523960 71946 524012 71952
rect 499856 71936 499908 71942
rect 499856 71878 499908 71884
rect 427728 71868 427780 71874
rect 427728 71810 427780 71816
rect 403624 71800 403676 71806
rect 403624 71742 403676 71748
rect 379520 71664 379572 71670
rect 379520 71606 379572 71612
rect 355600 71596 355652 71602
rect 355600 71538 355652 71544
rect 296076 71528 296128 71534
rect 296076 71470 296128 71476
rect 300952 71528 301004 71534
rect 300952 71470 301004 71476
rect 331496 71528 331548 71534
rect 331496 71470 331548 71476
rect 270592 3664 270644 3670
rect 270592 3606 270644 3612
rect 583392 3664 583444 3670
rect 583392 3606 583444 3612
rect 583404 480 583432 3606
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3606 667936 3662 667992
rect 2962 653540 3018 653576
rect 2962 653520 2964 653540
rect 2964 653520 3016 653540
rect 3016 653520 3018 653540
rect 2962 595992 3018 596048
rect 2962 538600 3018 538656
rect 2962 481072 3018 481128
rect 89166 700032 89222 700088
rect 24306 699896 24362 699952
rect 218978 700168 219034 700224
rect 3698 610408 3754 610464
rect 121734 585928 121790 585984
rect 3790 553016 3846 553072
rect 27250 581168 27306 581224
rect 24858 545536 24914 545592
rect 268290 547712 268346 547768
rect 24950 509904 25006 509960
rect 3882 495488 3938 495544
rect 24858 473048 24914 473104
rect 24950 402056 25006 402112
rect 24674 234640 24730 234696
rect 24766 199008 24822 199064
rect 24858 163376 24914 163432
rect 268842 511944 268898 512000
rect 269302 440680 269358 440736
rect 269302 405320 269358 405376
rect 270222 353776 270278 353832
rect 270038 348744 270094 348800
rect 269946 339904 270002 339960
rect 270130 339768 270186 339824
rect 269670 339632 269726 339688
rect 269854 335552 269910 335608
rect 270130 335552 270186 335608
rect 269394 329840 269450 329896
rect 237010 276156 237012 276176
rect 237012 276156 237064 276176
rect 237064 276156 237066 276176
rect 237010 276120 237066 276156
rect 247222 276156 247224 276176
rect 247224 276156 247276 276176
rect 247276 276156 247278 276176
rect 247222 276120 247278 276156
rect 27250 270816 27306 270872
rect 268382 237360 268438 237416
rect 268382 201728 268438 201784
rect 270406 345208 270462 345264
rect 270314 324400 270370 324456
rect 270590 353776 270646 353832
rect 270590 350784 270646 350840
rect 270498 320728 270554 320784
rect 270222 236988 270224 237008
rect 270224 236988 270276 237008
rect 270276 236988 270278 237008
rect 270222 236952 270278 236988
rect 270406 236952 270462 237008
rect 270130 216280 270186 216336
rect 270222 206080 270278 206136
rect 270222 195744 270278 195800
rect 270406 195744 270462 195800
rect 269946 185408 270002 185464
rect 270222 185408 270278 185464
rect 270222 175072 270278 175128
rect 270406 175072 270462 175128
rect 268566 166096 268622 166152
rect 270222 164736 270278 164792
rect 270406 164736 270462 164792
rect 270130 134000 270186 134056
rect 270130 132504 270186 132560
rect 267922 130464 267978 130520
rect 24950 128016 25006 128072
rect 267922 95104 267978 95160
rect 24950 92384 25006 92440
rect 269670 72120 269726 72176
rect 269854 72120 269910 72176
rect 270682 333648 270738 333704
rect 272338 381928 272394 381984
rect 272614 342388 272616 342408
rect 272616 342388 272668 342408
rect 272668 342388 272670 342408
rect 272614 342352 272670 342388
rect 272614 327528 272670 327584
rect 270774 317736 270830 317792
rect 494794 699896 494850 699952
rect 579894 697992 579950 698048
rect 579158 674600 579214 674656
rect 578790 627680 578846 627736
rect 307574 586492 307630 586528
rect 307574 586472 307576 586492
rect 307576 586472 307628 586492
rect 307628 586472 307630 586492
rect 341522 586472 341578 586528
rect 289450 586372 289452 586392
rect 289452 586372 289504 586392
rect 289504 586372 289506 586392
rect 289450 586336 289506 586372
rect 289450 586064 289506 586120
rect 298650 586064 298706 586120
rect 276386 510892 276388 510912
rect 276388 510892 276440 510912
rect 276440 510892 276442 510912
rect 276386 510856 276442 510892
rect 273902 382200 273958 382256
rect 283286 510856 283342 510912
rect 279698 359216 279754 359272
rect 280618 359216 280674 359272
rect 276754 354864 276810 354920
rect 297270 382064 297326 382120
rect 365442 586336 365498 586392
rect 413650 586200 413706 586256
rect 461674 586064 461730 586120
rect 315394 580660 315396 580680
rect 315396 580660 315448 580680
rect 315448 580660 315450 580680
rect 315394 580624 315450 580660
rect 314106 565120 314162 565176
rect 314198 559272 314254 559328
rect 303894 385600 303950 385656
rect 286966 354864 287022 354920
rect 289174 354864 289230 354920
rect 291198 354864 291254 354920
rect 293222 354864 293278 354920
rect 293590 354864 293646 354920
rect 300950 354864 301006 354920
rect 306930 354864 306986 354920
rect 311530 352008 311586 352064
rect 296534 316240 296590 316296
rect 275926 315560 275982 315616
rect 277674 313384 277730 313440
rect 281170 313248 281226 313304
rect 284022 313248 284078 313304
rect 279698 313112 279754 313168
rect 275650 312704 275706 312760
rect 276570 312704 276626 312760
rect 276662 273672 276718 273728
rect 276662 71984 276718 72040
rect 289818 276664 289874 276720
rect 293590 276664 293646 276720
rect 286230 133864 286286 133920
rect 298558 316240 298614 316296
rect 310886 316240 310942 316296
rect 306746 315560 306802 315616
rect 304538 315424 304594 315480
rect 303250 312704 303306 312760
rect 304538 312704 304594 312760
rect 306838 272176 306894 272232
rect 313554 339904 313610 339960
rect 313554 330928 313610 330984
rect 300950 72020 300952 72040
rect 300952 72020 301004 72040
rect 301004 72020 301006 72040
rect 300950 71984 301006 72020
rect 313738 345752 313794 345808
rect 313738 336504 313794 336560
rect 313646 327528 313702 327584
rect 315854 544876 315910 544912
rect 315854 544856 315856 544876
rect 315856 544856 315908 544876
rect 315908 544856 315910 544876
rect 314106 522552 314162 522608
rect 314474 522552 314530 522608
rect 315486 509496 315542 509552
rect 314382 504872 314438 504928
rect 314566 504872 314622 504928
rect 315486 473048 315542 473104
rect 314290 412156 314292 412176
rect 314292 412156 314344 412176
rect 314344 412156 314346 412176
rect 314290 412120 314346 412156
rect 314658 412120 314714 412176
rect 316222 402056 316278 402112
rect 314382 401920 314438 401976
rect 314658 401920 314714 401976
rect 379518 382200 379574 382256
rect 523958 382064 524014 382120
rect 548062 381928 548118 381984
rect 314106 370912 314162 370968
rect 314290 370912 314346 370968
rect 313922 348744 313978 348800
rect 314198 345752 314254 345808
rect 314106 336504 314162 336560
rect 313830 330928 313886 330984
rect 314382 348744 314438 348800
rect 578790 580760 578846 580816
rect 560850 547712 560906 547768
rect 578790 533840 578846 533896
rect 559378 512080 559434 512136
rect 560850 440680 560906 440736
rect 314934 333784 314990 333840
rect 560850 405320 560906 405376
rect 578790 392944 578846 393000
rect 560850 385600 560906 385656
rect 579894 651072 579950 651128
rect 579894 604152 579950 604208
rect 579894 557232 579950 557288
rect 579894 510312 579950 510368
rect 579250 486784 579306 486840
rect 579894 463392 579950 463448
rect 579342 439864 579398 439920
rect 579802 416472 579858 416528
rect 438030 275984 438086 276040
rect 315026 270272 315082 270328
rect 314290 234640 314346 234696
rect 560850 237360 560906 237416
rect 558918 201728 558974 201784
rect 315026 199008 315082 199064
rect 315026 163376 315082 163432
rect 559378 130464 559434 130520
rect 315026 92404 315082 92440
rect 315026 92384 315028 92404
rect 315028 92384 315080 92404
rect 315080 92384 315082 92404
rect 560850 95104 560906 95160
<< metal3 >>
rect 218973 700226 219039 700229
rect 310646 700226 310652 700228
rect 218973 700224 310652 700226
rect 218973 700168 218978 700224
rect 219034 700168 310652 700224
rect 218973 700166 310652 700168
rect 218973 700163 219039 700166
rect 310646 700164 310652 700166
rect 310716 700164 310722 700228
rect 89161 700090 89227 700093
rect 311014 700090 311020 700092
rect 89161 700088 311020 700090
rect 89161 700032 89166 700088
rect 89222 700032 311020 700088
rect 89161 700030 311020 700032
rect 89161 700027 89227 700030
rect 311014 700028 311020 700030
rect 311084 700028 311090 700092
rect 24301 699954 24367 699957
rect 310830 699954 310836 699956
rect 24301 699952 310836 699954
rect 24301 699896 24306 699952
rect 24362 699896 310836 699952
rect 24301 699894 310836 699896
rect 24301 699891 24367 699894
rect 310830 699892 310836 699894
rect 310900 699892 310906 699956
rect 311934 699892 311940 699956
rect 312004 699954 312010 699956
rect 494789 699954 494855 699957
rect 312004 699952 494855 699954
rect 312004 699896 494794 699952
rect 494850 699896 494855 699952
rect 312004 699894 494855 699896
rect 312004 699892 312010 699894
rect 494789 699891 494855 699894
rect 579889 698050 579955 698053
rect 583520 698050 584960 698140
rect 579889 698048 584960 698050
rect 579889 697992 579894 698048
rect 579950 697992 584960 698048
rect 579889 697990 584960 697992
rect 579889 697987 579955 697990
rect 583520 697900 584960 697990
rect -960 696540 480 696780
rect 583520 686204 584960 686444
rect -960 682124 480 682364
rect 579153 674658 579219 674661
rect 583520 674658 584960 674748
rect 579153 674656 584960 674658
rect 579153 674600 579158 674656
rect 579214 674600 584960 674656
rect 579153 674598 584960 674600
rect 579153 674595 579219 674598
rect 583520 674508 584960 674598
rect -960 667994 480 668084
rect 3601 667994 3667 667997
rect -960 667992 3667 667994
rect -960 667936 3606 667992
rect 3662 667936 3667 667992
rect -960 667934 3667 667936
rect -960 667844 480 667934
rect 3601 667931 3667 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 2957 653578 3023 653581
rect -960 653576 3023 653578
rect -960 653520 2962 653576
rect 3018 653520 3023 653576
rect -960 653518 3023 653520
rect -960 653428 480 653518
rect 2957 653515 3023 653518
rect 579889 651130 579955 651133
rect 583520 651130 584960 651220
rect 579889 651128 584960 651130
rect 579889 651072 579894 651128
rect 579950 651072 584960 651128
rect 579889 651070 584960 651072
rect 579889 651067 579955 651070
rect 583520 650980 584960 651070
rect 583520 639284 584960 639524
rect -960 639012 480 639252
rect 578785 627738 578851 627741
rect 583520 627738 584960 627828
rect 578785 627736 584960 627738
rect 578785 627680 578790 627736
rect 578846 627680 584960 627736
rect 578785 627678 584960 627680
rect 578785 627675 578851 627678
rect 583520 627588 584960 627678
rect -960 624732 480 624972
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 3693 610466 3759 610469
rect -960 610464 3759 610466
rect -960 610408 3698 610464
rect 3754 610408 3759 610464
rect -960 610406 3759 610408
rect -960 610316 480 610406
rect 3693 610403 3759 610406
rect 579889 604210 579955 604213
rect 583520 604210 584960 604300
rect 579889 604208 584960 604210
rect 579889 604152 579894 604208
rect 579950 604152 584960 604208
rect 579889 604150 584960 604152
rect 579889 604147 579955 604150
rect 583520 604060 584960 604150
rect -960 596050 480 596140
rect 2957 596050 3023 596053
rect -960 596048 3023 596050
rect -960 595992 2962 596048
rect 3018 595992 3023 596048
rect -960 595990 3023 595992
rect -960 595900 480 595990
rect 2957 595987 3023 595990
rect 583520 592364 584960 592604
rect 306598 586468 306604 586532
rect 306668 586530 306674 586532
rect 307569 586530 307635 586533
rect 341517 586530 341583 586533
rect 306668 586528 341583 586530
rect 306668 586472 307574 586528
rect 307630 586472 341522 586528
rect 341578 586472 341583 586528
rect 306668 586470 341583 586472
rect 306668 586468 306674 586470
rect 307569 586467 307635 586470
rect 341517 586467 341583 586470
rect 289445 586394 289511 586397
rect 365437 586394 365503 586397
rect 289445 586392 365503 586394
rect 289445 586336 289450 586392
rect 289506 586336 365442 586392
rect 365498 586336 365503 586392
rect 289445 586334 365503 586336
rect 289445 586331 289511 586334
rect 365437 586331 365503 586334
rect 289670 586196 289676 586260
rect 289740 586258 289746 586260
rect 413645 586258 413711 586261
rect 289740 586256 413711 586258
rect 289740 586200 413650 586256
rect 413706 586200 413711 586256
rect 289740 586198 413711 586200
rect 289740 586196 289746 586198
rect 413645 586195 413711 586198
rect 289445 586124 289511 586125
rect 298645 586124 298711 586125
rect 289445 586120 289492 586124
rect 289556 586122 289562 586124
rect 298645 586122 298692 586124
rect 289445 586064 289450 586120
rect 289445 586060 289492 586064
rect 289556 586062 289602 586122
rect 298564 586120 298692 586122
rect 298756 586122 298762 586124
rect 461669 586122 461735 586125
rect 298756 586120 461735 586122
rect 298564 586064 298650 586120
rect 298756 586064 461674 586120
rect 461730 586064 461735 586120
rect 298564 586062 298692 586064
rect 289556 586060 289562 586062
rect 298645 586060 298692 586062
rect 298756 586062 461735 586064
rect 298756 586060 298762 586062
rect 289445 586059 289511 586060
rect 298645 586059 298711 586060
rect 461669 586059 461735 586062
rect 121729 585986 121795 585989
rect 311198 585986 311204 585988
rect 121729 585984 311204 585986
rect 121729 585928 121734 585984
rect 121790 585928 311204 585984
rect 121729 585926 311204 585928
rect 121729 585923 121795 585926
rect 311198 585924 311204 585926
rect 311268 585924 311274 585988
rect -960 581620 480 581860
rect 27245 581226 27311 581229
rect 27245 581224 27354 581226
rect 27245 581168 27250 581224
rect 27306 581168 27354 581224
rect 27245 581163 27354 581168
rect 27294 580584 27354 581163
rect 578785 580818 578851 580821
rect 583520 580818 584960 580908
rect 578785 580816 584960 580818
rect 578785 580760 578790 580816
rect 578846 580760 584960 580816
rect 578785 580758 584960 580760
rect 578785 580755 578851 580758
rect 315389 580682 315455 580685
rect 315389 580680 318994 580682
rect 315389 580624 315394 580680
rect 315450 580624 318994 580680
rect 583520 580668 584960 580758
rect 315389 580622 318994 580624
rect 315389 580619 315455 580622
rect 318934 580584 318994 580622
rect 583520 568836 584960 569076
rect -960 567204 480 567444
rect 314101 565180 314167 565181
rect 314101 565176 314148 565180
rect 314212 565178 314218 565180
rect 314101 565120 314106 565176
rect 314101 565116 314148 565120
rect 314212 565118 314258 565178
rect 314212 565116 314218 565118
rect 314101 565115 314167 565116
rect 314193 559332 314259 559333
rect 314142 559330 314148 559332
rect 314102 559270 314148 559330
rect 314212 559328 314259 559332
rect 314254 559272 314259 559328
rect 314142 559268 314148 559270
rect 314212 559268 314259 559272
rect 314193 559267 314259 559268
rect 579889 557290 579955 557293
rect 583520 557290 584960 557380
rect 579889 557288 584960 557290
rect 579889 557232 579894 557288
rect 579950 557232 584960 557288
rect 579889 557230 584960 557232
rect 579889 557227 579955 557230
rect 583520 557140 584960 557230
rect -960 553074 480 553164
rect 3785 553074 3851 553077
rect -960 553072 3851 553074
rect -960 553016 3790 553072
rect 3846 553016 3851 553072
rect -960 553014 3851 553016
rect -960 552924 480 553014
rect 3785 553011 3851 553014
rect 268285 547770 268351 547773
rect 560845 547770 560911 547773
rect 266862 547768 268351 547770
rect 266862 547712 268290 547768
rect 268346 547712 268351 547768
rect 266862 547710 268351 547712
rect 266862 547702 266922 547710
rect 268285 547707 268351 547710
rect 558870 547768 560911 547770
rect 558870 547712 560850 547768
rect 560906 547712 560911 547768
rect 558870 547710 560911 547712
rect 558870 547702 558930 547710
rect 560845 547707 560911 547710
rect 266524 547642 266922 547702
rect 558716 547642 558930 547702
rect 24853 545594 24919 545597
rect 24853 545592 26802 545594
rect 24853 545536 24858 545592
rect 24914 545536 26802 545592
rect 24853 545534 26802 545536
rect 24853 545531 24919 545534
rect 26742 544952 26802 545534
rect 583520 545444 584960 545684
rect 315849 544914 315915 544917
rect 318934 544914 318994 544952
rect 315849 544912 318994 544914
rect 315849 544856 315854 544912
rect 315910 544856 318994 544912
rect 315849 544854 318994 544856
rect 315849 544851 315915 544854
rect -960 538658 480 538748
rect 2957 538658 3023 538661
rect -960 538656 3023 538658
rect -960 538600 2962 538656
rect 3018 538600 3023 538656
rect -960 538598 3023 538600
rect -960 538508 480 538598
rect 2957 538595 3023 538598
rect 578785 533898 578851 533901
rect 583520 533898 584960 533988
rect 578785 533896 584960 533898
rect 578785 533840 578790 533896
rect 578846 533840 584960 533896
rect 578785 533838 584960 533840
rect 578785 533835 578851 533838
rect 583520 533748 584960 533838
rect -960 524092 480 524332
rect 314101 522610 314167 522613
rect 314469 522610 314535 522613
rect 314101 522608 314535 522610
rect 314101 522552 314106 522608
rect 314162 522552 314474 522608
rect 314530 522552 314535 522608
rect 314101 522550 314535 522552
rect 314101 522547 314167 522550
rect 314469 522547 314535 522550
rect 583520 521916 584960 522156
rect 559373 512138 559439 512141
rect 558870 512136 559439 512138
rect 558870 512080 559378 512136
rect 559434 512080 559439 512136
rect 558870 512078 559439 512080
rect 558870 512070 558930 512078
rect 559373 512075 559439 512078
rect 266524 512010 266922 512070
rect 558716 512010 558930 512070
rect 266862 512002 266922 512010
rect 268837 512002 268903 512005
rect 266862 512000 268903 512002
rect 266862 511944 268842 512000
rect 268898 511944 268903 512000
rect 266862 511942 268903 511944
rect 268837 511939 268903 511942
rect 276381 510916 276447 510917
rect 276381 510914 276428 510916
rect 276336 510912 276428 510914
rect 276492 510914 276498 510916
rect 283281 510914 283347 510917
rect 276492 510912 283347 510914
rect 276336 510856 276386 510912
rect 276492 510856 283286 510912
rect 283342 510856 283347 510912
rect 276336 510854 276428 510856
rect 276381 510852 276428 510854
rect 276492 510854 283347 510856
rect 276492 510852 276498 510854
rect 276381 510851 276447 510852
rect 283281 510851 283347 510854
rect 579889 510370 579955 510373
rect 583520 510370 584960 510460
rect 579889 510368 584960 510370
rect 579889 510312 579894 510368
rect 579950 510312 584960 510368
rect 579889 510310 584960 510312
rect 579889 510307 579955 510310
rect 583520 510220 584960 510310
rect -960 509812 480 510052
rect 24945 509962 25011 509965
rect 24945 509960 26802 509962
rect 24945 509904 24950 509960
rect 25006 509904 26802 509960
rect 24945 509902 26802 509904
rect 24945 509899 25011 509902
rect 26742 509320 26802 509902
rect 315481 509554 315547 509557
rect 315481 509552 318994 509554
rect 315481 509496 315486 509552
rect 315542 509496 318994 509552
rect 315481 509494 318994 509496
rect 315481 509491 315547 509494
rect 318934 509320 318994 509494
rect 314377 504930 314443 504933
rect 314561 504930 314627 504933
rect 314377 504928 314627 504930
rect 314377 504872 314382 504928
rect 314438 504872 314566 504928
rect 314622 504872 314627 504928
rect 314377 504870 314627 504872
rect 314377 504867 314443 504870
rect 314561 504867 314627 504870
rect 583520 498524 584960 498764
rect -960 495546 480 495636
rect 3877 495546 3943 495549
rect -960 495544 3943 495546
rect -960 495488 3882 495544
rect 3938 495488 3943 495544
rect -960 495486 3943 495488
rect -960 495396 480 495486
rect 3877 495483 3943 495486
rect 579245 486842 579311 486845
rect 583520 486842 584960 486932
rect 579245 486840 584960 486842
rect 579245 486784 579250 486840
rect 579306 486784 584960 486840
rect 579245 486782 584960 486784
rect 579245 486779 579311 486782
rect 583520 486692 584960 486782
rect -960 481130 480 481220
rect 2957 481130 3023 481133
rect -960 481128 3023 481130
rect -960 481072 2962 481128
rect 3018 481072 3023 481128
rect -960 481070 3023 481072
rect -960 480980 480 481070
rect 2957 481067 3023 481070
rect 583520 474996 584960 475236
rect 24853 473106 24919 473109
rect 26742 473106 26802 473688
rect 24853 473104 26802 473106
rect 24853 473048 24858 473104
rect 24914 473048 26802 473104
rect 24853 473046 26802 473048
rect 315481 473106 315547 473109
rect 318934 473106 318994 473688
rect 315481 473104 318994 473106
rect 315481 473048 315486 473104
rect 315542 473048 318994 473104
rect 315481 473046 318994 473048
rect 24853 473043 24919 473046
rect 315481 473043 315547 473046
rect -960 466700 480 466940
rect 579889 463450 579955 463453
rect 583520 463450 584960 463540
rect 579889 463448 584960 463450
rect 579889 463392 579894 463448
rect 579950 463392 584960 463448
rect 579889 463390 584960 463392
rect 579889 463387 579955 463390
rect 583520 463300 584960 463390
rect -960 452284 480 452524
rect 583520 451604 584960 451844
rect 266524 440746 266922 440806
rect 558716 440746 559298 440806
rect 266862 440738 266922 440746
rect 269297 440738 269363 440741
rect 266862 440736 269363 440738
rect 266862 440680 269302 440736
rect 269358 440680 269363 440736
rect 266862 440678 269363 440680
rect 559238 440738 559298 440746
rect 560845 440738 560911 440741
rect 559238 440736 560911 440738
rect 559238 440680 560850 440736
rect 560906 440680 560911 440736
rect 559238 440678 560911 440680
rect 269297 440675 269363 440678
rect 560845 440675 560911 440678
rect 579337 439922 579403 439925
rect 583520 439922 584960 440012
rect 579337 439920 584960 439922
rect 579337 439864 579342 439920
rect 579398 439864 584960 439920
rect 579337 439862 584960 439864
rect 579337 439859 579403 439862
rect 583520 439772 584960 439862
rect -960 437868 480 438108
rect 583520 428076 584960 428316
rect -960 423588 480 423828
rect 579797 416530 579863 416533
rect 583520 416530 584960 416620
rect 579797 416528 584960 416530
rect 579797 416472 579802 416528
rect 579858 416472 584960 416528
rect 579797 416470 584960 416472
rect 579797 416467 579863 416470
rect 583520 416380 584960 416470
rect 314285 412178 314351 412181
rect 314653 412178 314719 412181
rect 314285 412176 314719 412178
rect 314285 412120 314290 412176
rect 314346 412120 314658 412176
rect 314714 412120 314719 412176
rect 314285 412118 314719 412120
rect 314285 412115 314351 412118
rect 314653 412115 314719 412118
rect -960 409172 480 409412
rect 266524 405386 266922 405446
rect 558716 405386 559298 405446
rect 266862 405378 266922 405386
rect 269297 405378 269363 405381
rect 266862 405376 269363 405378
rect 266862 405320 269302 405376
rect 269358 405320 269363 405376
rect 266862 405318 269363 405320
rect 559238 405378 559298 405386
rect 560845 405378 560911 405381
rect 559238 405376 560911 405378
rect 559238 405320 560850 405376
rect 560906 405320 560911 405376
rect 559238 405318 560911 405320
rect 269297 405315 269363 405318
rect 560845 405315 560911 405318
rect 583520 404684 584960 404924
rect 24945 402114 25011 402117
rect 26742 402114 26802 402696
rect 24945 402112 26802 402114
rect 24945 402056 24950 402112
rect 25006 402056 26802 402112
rect 24945 402054 26802 402056
rect 316217 402114 316283 402117
rect 318934 402114 318994 402696
rect 316217 402112 318994 402114
rect 316217 402056 316222 402112
rect 316278 402056 318994 402112
rect 316217 402054 318994 402056
rect 24945 402051 25011 402054
rect 316217 402051 316283 402054
rect 314377 401978 314443 401981
rect 314653 401978 314719 401981
rect 314377 401976 314719 401978
rect 314377 401920 314382 401976
rect 314438 401920 314658 401976
rect 314714 401920 314719 401976
rect 314377 401918 314719 401920
rect 314377 401915 314443 401918
rect 314653 401915 314719 401918
rect -960 394892 480 395132
rect 578785 393002 578851 393005
rect 583520 393002 584960 393092
rect 578785 393000 584960 393002
rect 578785 392944 578790 393000
rect 578846 392944 584960 393000
rect 578785 392942 584960 392944
rect 578785 392939 578851 392942
rect 583520 392852 584960 392942
rect 303889 385658 303955 385661
rect 304574 385658 304580 385660
rect 303889 385656 304580 385658
rect 303889 385600 303894 385656
rect 303950 385600 304580 385656
rect 303889 385598 304580 385600
rect 303889 385595 303955 385598
rect 304574 385596 304580 385598
rect 304644 385658 304650 385660
rect 560845 385658 560911 385661
rect 304644 385656 560911 385658
rect 304644 385600 560850 385656
rect 560906 385600 560911 385656
rect 304644 385598 560911 385600
rect 304644 385596 304650 385598
rect 560845 385595 560911 385598
rect 273897 382258 273963 382261
rect 275134 382258 275140 382260
rect 273897 382256 275140 382258
rect 273897 382200 273902 382256
rect 273958 382200 275140 382256
rect 273897 382198 275140 382200
rect 273897 382195 273963 382198
rect 275134 382196 275140 382198
rect 275204 382258 275210 382260
rect 379513 382258 379579 382261
rect 275204 382256 379579 382258
rect 275204 382200 379518 382256
rect 379574 382200 379579 382256
rect 275204 382198 379579 382200
rect 275204 382196 275210 382198
rect 379513 382195 379579 382198
rect 297265 382124 297331 382125
rect 297214 382122 297220 382124
rect 297138 382062 297220 382122
rect 297284 382122 297331 382124
rect 523953 382122 524019 382125
rect 297284 382120 524019 382122
rect 297326 382064 523958 382120
rect 524014 382064 524019 382120
rect 297214 382060 297220 382062
rect 297284 382062 524019 382064
rect 297284 382060 297331 382062
rect 297265 382059 297331 382060
rect 523953 382059 524019 382062
rect 272333 381986 272399 381989
rect 274950 381986 274956 381988
rect 272333 381984 274956 381986
rect 272333 381928 272338 381984
rect 272394 381928 274956 381984
rect 272333 381926 274956 381928
rect 272333 381923 272399 381926
rect 274950 381924 274956 381926
rect 275020 381986 275026 381988
rect 548057 381986 548123 381989
rect 275020 381984 548123 381986
rect 275020 381928 548062 381984
rect 548118 381928 548123 381984
rect 275020 381926 548123 381928
rect 275020 381924 275026 381926
rect 548057 381923 548123 381926
rect 583520 381156 584960 381396
rect -960 380476 480 380716
rect 314101 370970 314167 370973
rect 314285 370970 314351 370973
rect 314101 370968 314351 370970
rect 314101 370912 314106 370968
rect 314162 370912 314290 370968
rect 314346 370912 314351 370968
rect 314101 370910 314351 370912
rect 314101 370907 314167 370910
rect 314285 370907 314351 370910
rect 583520 369460 584960 369700
rect -960 366060 480 366300
rect 276606 359212 276612 359276
rect 276676 359274 276682 359276
rect 279693 359274 279759 359277
rect 280613 359274 280679 359277
rect 276676 359272 280679 359274
rect 276676 359216 279698 359272
rect 279754 359216 280618 359272
rect 280674 359216 280679 359272
rect 276676 359214 280679 359216
rect 276676 359212 276682 359214
rect 279693 359211 279759 359214
rect 280613 359211 280679 359214
rect 583520 357764 584960 358004
rect 275870 354860 275876 354924
rect 275940 354922 275946 354924
rect 276749 354922 276815 354925
rect 275940 354920 276815 354922
rect 275940 354864 276754 354920
rect 276810 354864 276815 354920
rect 275940 354862 276815 354864
rect 275940 354860 275946 354862
rect 276749 354859 276815 354862
rect 286961 354922 287027 354925
rect 287830 354922 287836 354924
rect 286961 354920 287836 354922
rect 286961 354864 286966 354920
rect 287022 354864 287836 354920
rect 286961 354862 287836 354864
rect 286961 354859 287027 354862
rect 287830 354860 287836 354862
rect 287900 354860 287906 354924
rect 289169 354922 289235 354925
rect 289854 354922 289860 354924
rect 289169 354920 289860 354922
rect 289169 354864 289174 354920
rect 289230 354864 289860 354920
rect 289169 354862 289860 354864
rect 289169 354859 289235 354862
rect 289854 354860 289860 354862
rect 289924 354860 289930 354924
rect 291193 354922 291259 354925
rect 291326 354922 291332 354924
rect 291193 354920 291332 354922
rect 291193 354864 291198 354920
rect 291254 354864 291332 354920
rect 291193 354862 291332 354864
rect 291193 354859 291259 354862
rect 291326 354860 291332 354862
rect 291396 354860 291402 354924
rect 293217 354922 293283 354925
rect 293585 354924 293651 354925
rect 300945 354924 301011 354925
rect 293534 354922 293540 354924
rect 293217 354920 293540 354922
rect 293604 354922 293651 354924
rect 293604 354920 293732 354922
rect 293217 354864 293222 354920
rect 293278 354864 293540 354920
rect 293646 354864 293732 354920
rect 293217 354862 293540 354864
rect 293217 354859 293283 354862
rect 293534 354860 293540 354862
rect 293604 354862 293732 354864
rect 293604 354860 293651 354862
rect 300894 354860 300900 354924
rect 300964 354922 301011 354924
rect 300964 354920 301056 354922
rect 301006 354864 301056 354920
rect 300964 354862 301056 354864
rect 300964 354860 301011 354862
rect 306414 354860 306420 354924
rect 306484 354922 306490 354924
rect 306925 354922 306991 354925
rect 306484 354920 306991 354922
rect 306484 354864 306930 354920
rect 306986 354864 306991 354920
rect 306484 354862 306991 354864
rect 306484 354860 306490 354862
rect 293585 354859 293651 354860
rect 300945 354859 301011 354860
rect 306925 354859 306991 354862
rect 270217 353834 270283 353837
rect 270585 353834 270651 353837
rect 272014 353834 272074 354348
rect 270217 353832 272074 353834
rect 270217 353776 270222 353832
rect 270278 353776 270590 353832
rect 270646 353776 272074 353832
rect 270217 353774 272074 353776
rect 270217 353771 270283 353774
rect 270585 353771 270651 353774
rect 311525 352066 311591 352069
rect 311525 352064 311634 352066
rect -960 351780 480 352020
rect 311525 352008 311530 352064
rect 311586 352008 311634 352064
rect 311525 352003 311634 352008
rect 311574 351628 311634 352003
rect 270585 350842 270651 350845
rect 272014 350842 272074 351356
rect 270585 350840 272074 350842
rect 270585 350784 270590 350840
rect 270646 350784 272074 350840
rect 270585 350782 272074 350784
rect 270585 350779 270651 350782
rect 270033 348802 270099 348805
rect 313917 348802 313983 348805
rect 314377 348802 314443 348805
rect 270033 348800 272074 348802
rect 270033 348744 270038 348800
rect 270094 348744 272074 348800
rect 270033 348742 272074 348744
rect 270033 348739 270099 348742
rect 272014 348364 272074 348742
rect 311942 348800 314443 348802
rect 311942 348744 313922 348800
rect 313978 348744 314382 348800
rect 314438 348744 314443 348800
rect 311942 348742 314443 348744
rect 311942 348636 312002 348742
rect 313917 348739 313983 348742
rect 314377 348739 314443 348742
rect 583520 345932 584960 346172
rect 313733 345810 313799 345813
rect 314193 345810 314259 345813
rect 311942 345808 314259 345810
rect 311942 345752 313738 345808
rect 313794 345752 314198 345808
rect 314254 345752 314259 345808
rect 311942 345750 314259 345752
rect 311942 345644 312002 345750
rect 313733 345747 313799 345750
rect 314193 345747 314259 345750
rect 270401 345266 270467 345269
rect 272014 345266 272074 345372
rect 270401 345264 272074 345266
rect 270401 345208 270406 345264
rect 270462 345208 272074 345264
rect 270401 345206 272074 345208
rect 270401 345203 270467 345206
rect 311566 343028 311572 343092
rect 311636 343028 311642 343092
rect 311574 342652 311634 343028
rect 272609 342410 272675 342413
rect 272566 342408 272675 342410
rect 272566 342352 272614 342408
rect 272670 342352 272675 342408
rect 272566 342347 272675 342352
rect 272566 342108 272626 342347
rect 269941 339960 270007 339965
rect 313549 339962 313615 339965
rect 269941 339904 269946 339960
rect 270002 339904 270007 339960
rect 269941 339899 270007 339904
rect 311942 339960 313615 339962
rect 311942 339904 313554 339960
rect 313610 339904 313615 339960
rect 311942 339902 313615 339904
rect 269944 339826 270004 339899
rect 270125 339826 270191 339829
rect 269944 339824 270191 339826
rect 269944 339768 270130 339824
rect 270186 339768 270191 339824
rect 269944 339766 270191 339768
rect 270125 339763 270191 339766
rect 269665 339690 269731 339693
rect 269665 339688 272074 339690
rect 269665 339632 269670 339688
rect 269726 339632 272074 339688
rect 311942 339660 312002 339902
rect 313549 339899 313615 339902
rect 269665 339630 272074 339632
rect 269665 339627 269731 339630
rect 272014 339116 272074 339630
rect -960 337364 480 337604
rect 313733 336562 313799 336565
rect 314101 336562 314167 336565
rect 311942 336560 314167 336562
rect 311942 336504 313738 336560
rect 313794 336504 314106 336560
rect 314162 336504 314167 336560
rect 311942 336502 314167 336504
rect 311942 336396 312002 336502
rect 313733 336499 313799 336502
rect 314101 336499 314167 336502
rect 269849 335610 269915 335613
rect 270125 335610 270191 335613
rect 272014 335610 272074 336124
rect 269849 335608 272074 335610
rect 269849 335552 269854 335608
rect 269910 335552 270130 335608
rect 270186 335552 272074 335608
rect 269849 335550 272074 335552
rect 269849 335547 269915 335550
rect 270125 335547 270191 335550
rect 583520 334236 584960 334476
rect 314929 333842 314995 333845
rect 311942 333840 314995 333842
rect 311942 333784 314934 333840
rect 314990 333784 314995 333840
rect 311942 333782 314995 333784
rect 270677 333706 270743 333709
rect 270677 333704 272074 333706
rect 270677 333648 270682 333704
rect 270738 333648 272074 333704
rect 270677 333646 272074 333648
rect 270677 333643 270743 333646
rect 272014 333132 272074 333646
rect 311942 333404 312002 333782
rect 314929 333779 314995 333782
rect 313549 330986 313615 330989
rect 313825 330986 313891 330989
rect 311942 330984 313891 330986
rect 311942 330928 313554 330984
rect 313610 330928 313830 330984
rect 313886 330928 313891 330984
rect 311942 330926 313891 330928
rect 311942 330412 312002 330926
rect 313549 330923 313615 330926
rect 313825 330923 313891 330926
rect 269389 329898 269455 329901
rect 272014 329898 272074 330140
rect 269389 329896 272074 329898
rect 269389 329840 269394 329896
rect 269450 329840 272074 329896
rect 269389 329838 272074 329840
rect 269389 329835 269455 329838
rect 272609 327586 272675 327589
rect 313641 327586 313707 327589
rect 272566 327584 272675 327586
rect 272566 327528 272614 327584
rect 272670 327528 272675 327584
rect 272566 327523 272675 327528
rect 311942 327584 313707 327586
rect 311942 327528 313646 327584
rect 313702 327528 313707 327584
rect 311942 327526 313707 327528
rect 272566 327148 272626 327523
rect 311942 327420 312002 327526
rect 313641 327523 313707 327526
rect 311566 324668 311572 324732
rect 311636 324668 311642 324732
rect 270309 324458 270375 324461
rect 270309 324456 272074 324458
rect 270309 324400 270314 324456
rect 270370 324400 272074 324456
rect 311574 324428 311634 324668
rect 270309 324398 272074 324400
rect 270309 324395 270375 324398
rect 272014 323884 272074 324398
rect -960 322948 480 323188
rect 583520 322540 584960 322780
rect 311566 321948 311572 322012
rect 311636 321948 311642 322012
rect 311574 321436 311634 321948
rect 270493 320786 270559 320789
rect 272014 320786 272074 320892
rect 270493 320784 272074 320786
rect 270493 320728 270498 320784
rect 270554 320728 272074 320784
rect 270493 320726 272074 320728
rect 270493 320723 270559 320726
rect 311566 318548 311572 318612
rect 311636 318548 311642 318612
rect 311574 318172 311634 318548
rect 270769 317794 270835 317797
rect 272014 317794 272074 317900
rect 270769 317792 272074 317794
rect 270769 317736 270774 317792
rect 270830 317736 272074 317792
rect 270769 317734 272074 317736
rect 270769 317731 270835 317734
rect 296529 316298 296595 316301
rect 297214 316298 297220 316300
rect 296529 316296 297220 316298
rect 296529 316240 296534 316296
rect 296590 316240 297220 316296
rect 296529 316238 297220 316240
rect 296529 316235 296595 316238
rect 297214 316236 297220 316238
rect 297284 316236 297290 316300
rect 298553 316298 298619 316301
rect 298686 316298 298692 316300
rect 298553 316296 298692 316298
rect 298553 316240 298558 316296
rect 298614 316240 298692 316296
rect 298553 316238 298692 316240
rect 298553 316235 298619 316238
rect 298686 316236 298692 316238
rect 298756 316236 298762 316300
rect 310881 316298 310947 316301
rect 311934 316298 311940 316300
rect 310881 316296 311940 316298
rect 310881 316240 310886 316296
rect 310942 316240 311940 316296
rect 310881 316238 311940 316240
rect 310881 316235 310947 316238
rect 311934 316236 311940 316238
rect 312004 316236 312010 316300
rect 275921 315618 275987 315621
rect 276422 315618 276428 315620
rect 275921 315616 276428 315618
rect 275921 315560 275926 315616
rect 275982 315560 276428 315616
rect 275921 315558 276428 315560
rect 275921 315555 275987 315558
rect 276422 315556 276428 315558
rect 276492 315556 276498 315620
rect 306598 315556 306604 315620
rect 306668 315618 306674 315620
rect 306741 315618 306807 315621
rect 306668 315616 306807 315618
rect 306668 315560 306746 315616
rect 306802 315560 306807 315616
rect 306668 315558 306807 315560
rect 306668 315556 306674 315558
rect 306741 315555 306807 315558
rect 304533 315484 304599 315485
rect 304533 315480 304580 315484
rect 304644 315482 304650 315484
rect 304533 315424 304538 315480
rect 304533 315420 304580 315424
rect 304644 315422 304690 315482
rect 304644 315420 304650 315422
rect 304533 315419 304599 315420
rect 277669 313442 277735 313445
rect 289670 313442 289676 313444
rect 277669 313440 289676 313442
rect 277669 313384 277674 313440
rect 277730 313384 289676 313440
rect 277669 313382 289676 313384
rect 277669 313379 277735 313382
rect 289670 313380 289676 313382
rect 289740 313380 289746 313444
rect 275134 313244 275140 313308
rect 275204 313306 275210 313308
rect 281165 313306 281231 313309
rect 275204 313304 281231 313306
rect 275204 313248 281170 313304
rect 281226 313248 281231 313304
rect 275204 313246 281231 313248
rect 275204 313244 275210 313246
rect 281165 313243 281231 313246
rect 284017 313306 284083 313309
rect 289486 313306 289492 313308
rect 284017 313304 289492 313306
rect 284017 313248 284022 313304
rect 284078 313248 289492 313304
rect 284017 313246 289492 313248
rect 284017 313243 284083 313246
rect 289486 313244 289492 313246
rect 289556 313244 289562 313308
rect 274950 313108 274956 313172
rect 275020 313170 275026 313172
rect 279693 313170 279759 313173
rect 275020 313168 279759 313170
rect 275020 313112 279698 313168
rect 279754 313112 279759 313168
rect 275020 313110 279759 313112
rect 275020 313108 275026 313110
rect 279693 313107 279759 313110
rect 275645 312762 275711 312765
rect 276565 312762 276631 312765
rect 275645 312760 276631 312762
rect 275645 312704 275650 312760
rect 275706 312704 276570 312760
rect 276626 312704 276631 312760
rect 275645 312702 276631 312704
rect 275645 312699 275711 312702
rect 276565 312699 276631 312702
rect 303245 312762 303311 312765
rect 304533 312762 304599 312765
rect 303245 312760 304599 312762
rect 303245 312704 303250 312760
rect 303306 312704 304538 312760
rect 304594 312704 304599 312760
rect 303245 312702 304599 312704
rect 303245 312699 303311 312702
rect 304533 312699 304599 312702
rect 583520 310708 584960 310948
rect -960 308668 480 308908
rect 583520 299012 584960 299252
rect -960 294252 480 294492
rect 583520 287316 584960 287556
rect -960 279972 480 280212
rect 289813 276724 289879 276725
rect 293585 276724 293651 276725
rect 289813 276720 289860 276724
rect 289924 276722 289930 276724
rect 293534 276722 293540 276724
rect 289813 276664 289818 276720
rect 289813 276660 289860 276664
rect 289924 276662 289970 276722
rect 293494 276662 293540 276722
rect 293604 276720 293651 276724
rect 293646 276664 293651 276720
rect 289924 276660 289930 276662
rect 293534 276660 293540 276662
rect 293604 276660 293651 276664
rect 289813 276659 289879 276660
rect 293585 276659 293651 276660
rect 237005 276178 237071 276181
rect 247217 276178 247283 276181
rect 237005 276176 247283 276178
rect 237005 276120 237010 276176
rect 237066 276120 247222 276176
rect 247278 276120 247283 276176
rect 237005 276118 247283 276120
rect 237005 276115 237071 276118
rect 247217 276115 247283 276118
rect 291326 275980 291332 276044
rect 291396 276042 291402 276044
rect 438025 276042 438091 276045
rect 291396 276040 438091 276042
rect 291396 275984 438030 276040
rect 438086 275984 438091 276040
rect 291396 275982 438091 275984
rect 291396 275980 291402 275982
rect 438025 275979 438091 275982
rect 583520 275620 584960 275860
rect 275870 273668 275876 273732
rect 275940 273730 275946 273732
rect 276657 273730 276723 273733
rect 275940 273728 276723 273730
rect 275940 273672 276662 273728
rect 276718 273672 276723 273728
rect 275940 273670 276723 273672
rect 275940 273668 275946 273670
rect 276657 273667 276723 273670
rect 306414 272172 306420 272236
rect 306484 272234 306490 272236
rect 306833 272234 306899 272237
rect 306484 272232 306899 272234
rect 306484 272176 306838 272232
rect 306894 272176 306899 272232
rect 306484 272174 306899 272176
rect 306484 272172 306490 272174
rect 306833 272171 306899 272174
rect 27245 270874 27311 270877
rect 27245 270872 27354 270874
rect 27245 270816 27250 270872
rect 27306 270816 27354 270872
rect 27245 270811 27354 270816
rect 27294 270300 27354 270811
rect 315021 270330 315087 270333
rect 315021 270328 318964 270330
rect 315021 270272 315026 270328
rect 315082 270272 318964 270328
rect 315021 270270 318964 270272
rect 315021 270267 315087 270270
rect -960 265556 480 265796
rect 583520 263788 584960 264028
rect 583520 252092 584960 252332
rect -960 251140 480 251380
rect 583520 240396 584960 240636
rect 268377 237418 268443 237421
rect 560845 237418 560911 237421
rect 266524 237416 268443 237418
rect 266524 237360 268382 237416
rect 268438 237360 268443 237416
rect 266524 237358 268443 237360
rect 558716 237416 560911 237418
rect 558716 237360 560850 237416
rect 560906 237360 560911 237416
rect 558716 237358 560911 237360
rect 268377 237355 268443 237358
rect 560845 237355 560911 237358
rect -960 236860 480 237100
rect 270217 237010 270283 237013
rect 270401 237010 270467 237013
rect 270217 237008 270467 237010
rect 270217 236952 270222 237008
rect 270278 236952 270406 237008
rect 270462 236952 270467 237008
rect 270217 236950 270467 236952
rect 270217 236947 270283 236950
rect 270401 236947 270467 236950
rect 24669 234698 24735 234701
rect 314285 234698 314351 234701
rect 24669 234696 26772 234698
rect 24669 234640 24674 234696
rect 24730 234640 26772 234696
rect 24669 234638 26772 234640
rect 314285 234696 318964 234698
rect 314285 234640 314290 234696
rect 314346 234640 318964 234696
rect 314285 234638 318964 234640
rect 24669 234635 24735 234638
rect 314285 234635 314351 234638
rect 583520 228700 584960 228940
rect -960 222444 480 222684
rect 583520 216868 584960 217108
rect 270125 216340 270191 216341
rect 270125 216336 270172 216340
rect 270236 216338 270242 216340
rect 270125 216280 270130 216336
rect 270125 216276 270172 216280
rect 270236 216278 270282 216338
rect 270236 216276 270242 216278
rect 270125 216275 270191 216276
rect -960 208028 480 208268
rect 270217 206140 270283 206141
rect 270166 206138 270172 206140
rect 270126 206078 270172 206138
rect 270236 206136 270283 206140
rect 270278 206080 270283 206136
rect 270166 206076 270172 206078
rect 270236 206076 270283 206080
rect 270217 206075 270283 206076
rect 583520 205172 584960 205412
rect 268377 201786 268443 201789
rect 558913 201786 558979 201789
rect 266524 201784 268443 201786
rect 266524 201728 268382 201784
rect 268438 201728 268443 201784
rect 266524 201726 268443 201728
rect 558716 201784 558979 201786
rect 558716 201728 558918 201784
rect 558974 201728 558979 201784
rect 558716 201726 558979 201728
rect 268377 201723 268443 201726
rect 558913 201723 558979 201726
rect 24761 199066 24827 199069
rect 315021 199066 315087 199069
rect 24761 199064 26772 199066
rect 24761 199008 24766 199064
rect 24822 199008 26772 199064
rect 24761 199006 26772 199008
rect 315021 199064 318964 199066
rect 315021 199008 315026 199064
rect 315082 199008 318964 199064
rect 315021 199006 318964 199008
rect 24761 199003 24827 199006
rect 315021 199003 315087 199006
rect 270217 195802 270283 195805
rect 270401 195802 270467 195805
rect 270217 195800 270467 195802
rect 270217 195744 270222 195800
rect 270278 195744 270406 195800
rect 270462 195744 270467 195800
rect 270217 195742 270467 195744
rect 270217 195739 270283 195742
rect 270401 195739 270467 195742
rect -960 193748 480 193988
rect 583520 193476 584960 193716
rect 269941 185466 270007 185469
rect 270217 185466 270283 185469
rect 269941 185464 270283 185466
rect 269941 185408 269946 185464
rect 270002 185408 270222 185464
rect 270278 185408 270283 185464
rect 269941 185406 270283 185408
rect 269941 185403 270007 185406
rect 270217 185403 270283 185406
rect 583520 181780 584960 182020
rect -960 179332 480 179572
rect 270217 175130 270283 175133
rect 270401 175130 270467 175133
rect 270217 175128 270467 175130
rect 270217 175072 270222 175128
rect 270278 175072 270406 175128
rect 270462 175072 270467 175128
rect 270217 175070 270467 175072
rect 270217 175067 270283 175070
rect 270401 175067 270467 175070
rect 583520 169948 584960 170188
rect 268561 166154 268627 166157
rect 266524 166152 268627 166154
rect 266524 166096 268566 166152
rect 268622 166096 268627 166152
rect 266524 166094 268627 166096
rect 268561 166091 268627 166094
rect -960 164916 480 165156
rect 270217 164794 270283 164797
rect 270401 164794 270467 164797
rect 270217 164792 270467 164794
rect 270217 164736 270222 164792
rect 270278 164736 270406 164792
rect 270462 164736 270467 164792
rect 270217 164734 270467 164736
rect 270217 164731 270283 164734
rect 270401 164731 270467 164734
rect 24853 163434 24919 163437
rect 315021 163434 315087 163437
rect 24853 163432 26772 163434
rect 24853 163376 24858 163432
rect 24914 163376 26772 163432
rect 24853 163374 26772 163376
rect 315021 163432 318964 163434
rect 315021 163376 315026 163432
rect 315082 163376 318964 163432
rect 315021 163374 318964 163376
rect 24853 163371 24919 163374
rect 315021 163371 315087 163374
rect 583520 158252 584960 158492
rect -960 150636 480 150876
rect 583520 146556 584960 146796
rect -960 136220 480 136460
rect 583520 134724 584960 134964
rect 270125 134060 270191 134061
rect 270125 134056 270172 134060
rect 270236 134058 270242 134060
rect 270125 134000 270130 134056
rect 270125 133996 270172 134000
rect 270236 133998 270282 134058
rect 270236 133996 270242 133998
rect 270125 133995 270191 133996
rect 286225 133922 286291 133925
rect 287830 133922 287836 133924
rect 286225 133920 287836 133922
rect 286225 133864 286230 133920
rect 286286 133864 287836 133920
rect 286225 133862 287836 133864
rect 286225 133859 286291 133862
rect 287830 133860 287836 133862
rect 287900 133860 287906 133924
rect 270125 132564 270191 132565
rect 270125 132560 270172 132564
rect 270236 132562 270242 132564
rect 270125 132504 270130 132560
rect 270125 132500 270172 132504
rect 270236 132502 270282 132562
rect 270236 132500 270242 132502
rect 270125 132499 270191 132500
rect 267917 130522 267983 130525
rect 559373 130522 559439 130525
rect 266524 130520 267983 130522
rect 266524 130464 267922 130520
rect 267978 130464 267983 130520
rect 266524 130462 267983 130464
rect 558716 130520 559439 130522
rect 558716 130464 559378 130520
rect 559434 130464 559439 130520
rect 558716 130462 559439 130464
rect 267917 130459 267983 130462
rect 559373 130459 559439 130462
rect 24945 128074 25011 128077
rect 24945 128072 26772 128074
rect 24945 128016 24950 128072
rect 25006 128016 26772 128072
rect 24945 128014 26772 128016
rect 24945 128011 25011 128014
rect 583520 123028 584960 123268
rect -960 121940 480 122180
rect 583520 111332 584960 111572
rect -960 107524 480 107764
rect 583520 99636 584960 99876
rect 267917 95162 267983 95165
rect 560845 95162 560911 95165
rect 266524 95160 267983 95162
rect 266524 95104 267922 95160
rect 267978 95104 267983 95160
rect 266524 95102 267983 95104
rect 558716 95160 560911 95162
rect 558716 95104 560850 95160
rect 560906 95104 560911 95160
rect 558716 95102 560911 95104
rect 267917 95099 267983 95102
rect 560845 95099 560911 95102
rect -960 93108 480 93348
rect 24945 92442 25011 92445
rect 315021 92442 315087 92445
rect 24945 92440 26772 92442
rect 24945 92384 24950 92440
rect 25006 92384 26772 92440
rect 24945 92382 26772 92384
rect 315021 92440 318964 92442
rect 315021 92384 315026 92440
rect 315082 92384 318964 92440
rect 315021 92382 318964 92384
rect 24945 92379 25011 92382
rect 315021 92379 315087 92382
rect 583520 87804 584960 88044
rect -960 78828 480 79068
rect 583520 76108 584960 76348
rect 269665 72178 269731 72181
rect 269849 72178 269915 72181
rect 269665 72176 269915 72178
rect 269665 72120 269670 72176
rect 269726 72120 269854 72176
rect 269910 72120 269915 72176
rect 269665 72118 269915 72120
rect 269665 72115 269731 72118
rect 269849 72115 269915 72118
rect 276657 72044 276723 72045
rect 300945 72044 301011 72045
rect 276606 72042 276612 72044
rect 276566 71982 276612 72042
rect 276676 72040 276723 72044
rect 300894 72042 300900 72044
rect 276718 71984 276723 72040
rect 276606 71980 276612 71982
rect 276676 71980 276723 71984
rect 300854 71982 300900 72042
rect 300964 72040 301011 72044
rect 301006 71984 301011 72040
rect 300894 71980 300900 71982
rect 300964 71980 301011 71984
rect 276657 71979 276723 71980
rect 300945 71979 301011 71980
rect -960 64412 480 64652
rect 583520 64412 584960 64652
rect 583520 52716 584960 52956
rect -960 49996 480 50236
rect 583520 40884 584960 41124
rect -960 35716 480 35956
rect 583520 29188 584960 29428
rect -960 21300 480 21540
rect 583520 17492 584960 17732
rect -960 7020 480 7260
rect 583520 5796 584960 6036
<< via3 >>
rect 310652 700164 310716 700228
rect 311020 700028 311084 700092
rect 310836 699892 310900 699956
rect 311940 699892 312004 699956
rect 306604 586468 306668 586532
rect 289676 586196 289740 586260
rect 289492 586120 289556 586124
rect 289492 586064 289506 586120
rect 289506 586064 289556 586120
rect 289492 586060 289556 586064
rect 298692 586120 298756 586124
rect 298692 586064 298706 586120
rect 298706 586064 298756 586120
rect 298692 586060 298756 586064
rect 311204 585924 311268 585988
rect 314148 565176 314212 565180
rect 314148 565120 314162 565176
rect 314162 565120 314212 565176
rect 314148 565116 314212 565120
rect 314148 559328 314212 559332
rect 314148 559272 314198 559328
rect 314198 559272 314212 559328
rect 314148 559268 314212 559272
rect 276428 510912 276492 510916
rect 276428 510856 276442 510912
rect 276442 510856 276492 510912
rect 276428 510852 276492 510856
rect 304580 385596 304644 385660
rect 275140 382196 275204 382260
rect 297220 382120 297284 382124
rect 297220 382064 297270 382120
rect 297270 382064 297284 382120
rect 297220 382060 297284 382064
rect 274956 381924 275020 381988
rect 276612 359212 276676 359276
rect 275876 354860 275940 354924
rect 287836 354860 287900 354924
rect 289860 354860 289924 354924
rect 291332 354860 291396 354924
rect 293540 354920 293604 354924
rect 293540 354864 293590 354920
rect 293590 354864 293604 354920
rect 293540 354860 293604 354864
rect 300900 354920 300964 354924
rect 300900 354864 300950 354920
rect 300950 354864 300964 354920
rect 300900 354860 300964 354864
rect 306420 354860 306484 354924
rect 311572 343028 311636 343092
rect 311572 324668 311636 324732
rect 311572 321948 311636 322012
rect 311572 318548 311636 318612
rect 297220 316236 297284 316300
rect 298692 316236 298756 316300
rect 311940 316236 312004 316300
rect 276428 315556 276492 315620
rect 306604 315556 306668 315620
rect 304580 315480 304644 315484
rect 304580 315424 304594 315480
rect 304594 315424 304644 315480
rect 304580 315420 304644 315424
rect 289676 313380 289740 313444
rect 275140 313244 275204 313308
rect 289492 313244 289556 313308
rect 274956 313108 275020 313172
rect 289860 276720 289924 276724
rect 289860 276664 289874 276720
rect 289874 276664 289924 276720
rect 289860 276660 289924 276664
rect 293540 276720 293604 276724
rect 293540 276664 293590 276720
rect 293590 276664 293604 276720
rect 293540 276660 293604 276664
rect 291332 275980 291396 276044
rect 275876 273668 275940 273732
rect 306420 272172 306484 272236
rect 270172 216336 270236 216340
rect 270172 216280 270186 216336
rect 270186 216280 270236 216336
rect 270172 216276 270236 216280
rect 270172 206136 270236 206140
rect 270172 206080 270222 206136
rect 270222 206080 270236 206136
rect 270172 206076 270236 206080
rect 270172 134056 270236 134060
rect 270172 134000 270186 134056
rect 270186 134000 270236 134056
rect 270172 133996 270236 134000
rect 287836 133860 287900 133924
rect 270172 132560 270236 132564
rect 270172 132504 270186 132560
rect 270186 132504 270236 132560
rect 270172 132500 270236 132504
rect 276612 72040 276676 72044
rect 276612 71984 276662 72040
rect 276662 71984 276676 72040
rect 276612 71980 276676 71984
rect 300900 72040 300964 72044
rect 300900 71984 300950 72040
rect 300950 71984 300964 72040
rect 300900 71980 300964 71984
<< metal4 >>
rect -8576 711418 -7976 711440
rect -8576 711182 -8394 711418
rect -8158 711182 -7976 711418
rect -8576 711098 -7976 711182
rect -8576 710862 -8394 711098
rect -8158 710862 -7976 711098
rect -8576 -6926 -7976 710862
rect 591900 711418 592500 711440
rect 591900 711182 592082 711418
rect 592318 711182 592500 711418
rect 591900 711098 592500 711182
rect 591900 710862 592082 711098
rect 592318 710862 592500 711098
rect -7636 710478 -7036 710500
rect -7636 710242 -7454 710478
rect -7218 710242 -7036 710478
rect -7636 710158 -7036 710242
rect -7636 709922 -7454 710158
rect -7218 709922 -7036 710158
rect -7636 -5986 -7036 709922
rect 590960 710478 591560 710500
rect 590960 710242 591142 710478
rect 591378 710242 591560 710478
rect 590960 710158 591560 710242
rect 590960 709922 591142 710158
rect 591378 709922 591560 710158
rect -6696 709538 -6096 709560
rect -6696 709302 -6514 709538
rect -6278 709302 -6096 709538
rect -6696 709218 -6096 709302
rect -6696 708982 -6514 709218
rect -6278 708982 -6096 709218
rect -6696 -5046 -6096 708982
rect 590020 709538 590620 709560
rect 590020 709302 590202 709538
rect 590438 709302 590620 709538
rect 590020 709218 590620 709302
rect 590020 708982 590202 709218
rect 590438 708982 590620 709218
rect -5756 708598 -5156 708620
rect -5756 708362 -5574 708598
rect -5338 708362 -5156 708598
rect -5756 708278 -5156 708362
rect -5756 708042 -5574 708278
rect -5338 708042 -5156 708278
rect -5756 -4106 -5156 708042
rect 589080 708598 589680 708620
rect 589080 708362 589262 708598
rect 589498 708362 589680 708598
rect 589080 708278 589680 708362
rect 589080 708042 589262 708278
rect 589498 708042 589680 708278
rect -4816 707658 -4216 707680
rect -4816 707422 -4634 707658
rect -4398 707422 -4216 707658
rect -4816 707338 -4216 707422
rect -4816 707102 -4634 707338
rect -4398 707102 -4216 707338
rect -4816 -3166 -4216 707102
rect 588140 707658 588740 707680
rect 588140 707422 588322 707658
rect 588558 707422 588740 707658
rect 588140 707338 588740 707422
rect 588140 707102 588322 707338
rect 588558 707102 588740 707338
rect -3876 706718 -3276 706740
rect -3876 706482 -3694 706718
rect -3458 706482 -3276 706718
rect -3876 706398 -3276 706482
rect -3876 706162 -3694 706398
rect -3458 706162 -3276 706398
rect -3876 -2226 -3276 706162
rect 587200 706718 587800 706740
rect 587200 706482 587382 706718
rect 587618 706482 587800 706718
rect 587200 706398 587800 706482
rect 587200 706162 587382 706398
rect 587618 706162 587800 706398
rect -2936 705778 -2336 705800
rect -2936 705542 -2754 705778
rect -2518 705542 -2336 705778
rect -2936 705458 -2336 705542
rect -2936 705222 -2754 705458
rect -2518 705222 -2336 705458
rect -2936 668454 -2336 705222
rect -2936 668218 -2754 668454
rect -2518 668218 -2336 668454
rect -2936 668134 -2336 668218
rect -2936 667898 -2754 668134
rect -2518 667898 -2336 668134
rect -2936 632454 -2336 667898
rect -2936 632218 -2754 632454
rect -2518 632218 -2336 632454
rect -2936 632134 -2336 632218
rect -2936 631898 -2754 632134
rect -2518 631898 -2336 632134
rect -2936 596454 -2336 631898
rect -2936 596218 -2754 596454
rect -2518 596218 -2336 596454
rect -2936 596134 -2336 596218
rect -2936 595898 -2754 596134
rect -2518 595898 -2336 596134
rect -2936 560454 -2336 595898
rect -2936 560218 -2754 560454
rect -2518 560218 -2336 560454
rect -2936 560134 -2336 560218
rect -2936 559898 -2754 560134
rect -2518 559898 -2336 560134
rect -2936 524454 -2336 559898
rect -2936 524218 -2754 524454
rect -2518 524218 -2336 524454
rect -2936 524134 -2336 524218
rect -2936 523898 -2754 524134
rect -2518 523898 -2336 524134
rect -2936 488454 -2336 523898
rect -2936 488218 -2754 488454
rect -2518 488218 -2336 488454
rect -2936 488134 -2336 488218
rect -2936 487898 -2754 488134
rect -2518 487898 -2336 488134
rect -2936 452454 -2336 487898
rect -2936 452218 -2754 452454
rect -2518 452218 -2336 452454
rect -2936 452134 -2336 452218
rect -2936 451898 -2754 452134
rect -2518 451898 -2336 452134
rect -2936 416454 -2336 451898
rect -2936 416218 -2754 416454
rect -2518 416218 -2336 416454
rect -2936 416134 -2336 416218
rect -2936 415898 -2754 416134
rect -2518 415898 -2336 416134
rect -2936 380454 -2336 415898
rect -2936 380218 -2754 380454
rect -2518 380218 -2336 380454
rect -2936 380134 -2336 380218
rect -2936 379898 -2754 380134
rect -2518 379898 -2336 380134
rect -2936 344454 -2336 379898
rect -2936 344218 -2754 344454
rect -2518 344218 -2336 344454
rect -2936 344134 -2336 344218
rect -2936 343898 -2754 344134
rect -2518 343898 -2336 344134
rect -2936 308454 -2336 343898
rect -2936 308218 -2754 308454
rect -2518 308218 -2336 308454
rect -2936 308134 -2336 308218
rect -2936 307898 -2754 308134
rect -2518 307898 -2336 308134
rect -2936 272454 -2336 307898
rect -2936 272218 -2754 272454
rect -2518 272218 -2336 272454
rect -2936 272134 -2336 272218
rect -2936 271898 -2754 272134
rect -2518 271898 -2336 272134
rect -2936 236454 -2336 271898
rect -2936 236218 -2754 236454
rect -2518 236218 -2336 236454
rect -2936 236134 -2336 236218
rect -2936 235898 -2754 236134
rect -2518 235898 -2336 236134
rect -2936 200454 -2336 235898
rect -2936 200218 -2754 200454
rect -2518 200218 -2336 200454
rect -2936 200134 -2336 200218
rect -2936 199898 -2754 200134
rect -2518 199898 -2336 200134
rect -2936 164454 -2336 199898
rect -2936 164218 -2754 164454
rect -2518 164218 -2336 164454
rect -2936 164134 -2336 164218
rect -2936 163898 -2754 164134
rect -2518 163898 -2336 164134
rect -2936 128454 -2336 163898
rect -2936 128218 -2754 128454
rect -2518 128218 -2336 128454
rect -2936 128134 -2336 128218
rect -2936 127898 -2754 128134
rect -2518 127898 -2336 128134
rect -2936 92454 -2336 127898
rect -2936 92218 -2754 92454
rect -2518 92218 -2336 92454
rect -2936 92134 -2336 92218
rect -2936 91898 -2754 92134
rect -2518 91898 -2336 92134
rect -2936 56454 -2336 91898
rect -2936 56218 -2754 56454
rect -2518 56218 -2336 56454
rect -2936 56134 -2336 56218
rect -2936 55898 -2754 56134
rect -2518 55898 -2336 56134
rect -2936 20454 -2336 55898
rect -2936 20218 -2754 20454
rect -2518 20218 -2336 20454
rect -2936 20134 -2336 20218
rect -2936 19898 -2754 20134
rect -2518 19898 -2336 20134
rect -2936 -1286 -2336 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705800
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2936 -1522 -2754 -1286
rect -2518 -1522 -2336 -1286
rect -2936 -1606 -2336 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 -2336 -1606
rect -2936 -1864 -2336 -1842
rect 804 -1864 1404 -902
rect 18804 705778 19404 705800
rect 18804 705542 18986 705778
rect 19222 705542 19404 705778
rect 18804 705458 19404 705542
rect 18804 705222 18986 705458
rect 19222 705222 19404 705458
rect 18804 668454 19404 705222
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 36804 704838 37404 705800
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 584916 37404 613898
rect 54804 705778 55404 705800
rect 54804 705542 54986 705778
rect 55222 705542 55404 705778
rect 54804 705458 55404 705542
rect 54804 705222 54986 705458
rect 55222 705222 55404 705458
rect 54804 668454 55404 705222
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 584916 55404 595898
rect 72804 704838 73404 705800
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 614454 73404 649898
rect 72804 614218 72986 614454
rect 73222 614218 73404 614454
rect 72804 614134 73404 614218
rect 72804 613898 72986 614134
rect 73222 613898 73404 614134
rect 72804 584916 73404 613898
rect 90804 705778 91404 705800
rect 90804 705542 90986 705778
rect 91222 705542 91404 705778
rect 90804 705458 91404 705542
rect 90804 705222 90986 705458
rect 91222 705222 91404 705458
rect 90804 668454 91404 705222
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 632454 91404 667898
rect 90804 632218 90986 632454
rect 91222 632218 91404 632454
rect 90804 632134 91404 632218
rect 90804 631898 90986 632134
rect 91222 631898 91404 632134
rect 90804 596454 91404 631898
rect 90804 596218 90986 596454
rect 91222 596218 91404 596454
rect 90804 596134 91404 596218
rect 90804 595898 90986 596134
rect 91222 595898 91404 596134
rect 90804 584916 91404 595898
rect 108804 704838 109404 705800
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 650454 109404 685898
rect 108804 650218 108986 650454
rect 109222 650218 109404 650454
rect 108804 650134 109404 650218
rect 108804 649898 108986 650134
rect 109222 649898 109404 650134
rect 108804 614454 109404 649898
rect 108804 614218 108986 614454
rect 109222 614218 109404 614454
rect 108804 614134 109404 614218
rect 108804 613898 108986 614134
rect 109222 613898 109404 614134
rect 108804 584916 109404 613898
rect 126804 705778 127404 705800
rect 126804 705542 126986 705778
rect 127222 705542 127404 705778
rect 126804 705458 127404 705542
rect 126804 705222 126986 705458
rect 127222 705222 127404 705458
rect 126804 668454 127404 705222
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 632454 127404 667898
rect 126804 632218 126986 632454
rect 127222 632218 127404 632454
rect 126804 632134 127404 632218
rect 126804 631898 126986 632134
rect 127222 631898 127404 632134
rect 126804 596454 127404 631898
rect 126804 596218 126986 596454
rect 127222 596218 127404 596454
rect 126804 596134 127404 596218
rect 126804 595898 126986 596134
rect 127222 595898 127404 596134
rect 126804 584916 127404 595898
rect 144804 704838 145404 705800
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 144804 584916 145404 613898
rect 162804 705778 163404 705800
rect 162804 705542 162986 705778
rect 163222 705542 163404 705778
rect 162804 705458 163404 705542
rect 162804 705222 162986 705458
rect 163222 705222 163404 705458
rect 162804 668454 163404 705222
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 162804 584916 163404 595898
rect 180804 704838 181404 705800
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 584916 181404 613898
rect 198804 705778 199404 705800
rect 198804 705542 198986 705778
rect 199222 705542 199404 705778
rect 198804 705458 199404 705542
rect 198804 705222 198986 705458
rect 199222 705222 199404 705458
rect 198804 668454 199404 705222
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 632454 199404 667898
rect 198804 632218 198986 632454
rect 199222 632218 199404 632454
rect 198804 632134 199404 632218
rect 198804 631898 198986 632134
rect 199222 631898 199404 632134
rect 198804 596454 199404 631898
rect 198804 596218 198986 596454
rect 199222 596218 199404 596454
rect 198804 596134 199404 596218
rect 198804 595898 198986 596134
rect 199222 595898 199404 596134
rect 198804 584916 199404 595898
rect 216804 704838 217404 705800
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 650454 217404 685898
rect 216804 650218 216986 650454
rect 217222 650218 217404 650454
rect 216804 650134 217404 650218
rect 216804 649898 216986 650134
rect 217222 649898 217404 650134
rect 216804 614454 217404 649898
rect 216804 614218 216986 614454
rect 217222 614218 217404 614454
rect 216804 614134 217404 614218
rect 216804 613898 216986 614134
rect 217222 613898 217404 614134
rect 216804 584916 217404 613898
rect 234804 705778 235404 705800
rect 234804 705542 234986 705778
rect 235222 705542 235404 705778
rect 234804 705458 235404 705542
rect 234804 705222 234986 705458
rect 235222 705222 235404 705458
rect 234804 668454 235404 705222
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 632454 235404 667898
rect 234804 632218 234986 632454
rect 235222 632218 235404 632454
rect 234804 632134 235404 632218
rect 234804 631898 234986 632134
rect 235222 631898 235404 632134
rect 234804 596454 235404 631898
rect 234804 596218 234986 596454
rect 235222 596218 235404 596454
rect 234804 596134 235404 596218
rect 234804 595898 234986 596134
rect 235222 595898 235404 596134
rect 234804 584916 235404 595898
rect 252804 704838 253404 705800
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 650454 253404 685898
rect 252804 650218 252986 650454
rect 253222 650218 253404 650454
rect 252804 650134 253404 650218
rect 252804 649898 252986 650134
rect 253222 649898 253404 650134
rect 252804 614454 253404 649898
rect 252804 614218 252986 614454
rect 253222 614218 253404 614454
rect 252804 614134 253404 614218
rect 252804 613898 252986 614134
rect 253222 613898 253404 614134
rect 252804 584916 253404 613898
rect 270804 705778 271404 705800
rect 270804 705542 270986 705778
rect 271222 705542 271404 705778
rect 270804 705458 271404 705542
rect 270804 705222 270986 705458
rect 271222 705222 271404 705458
rect 270804 668454 271404 705222
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 270804 596454 271404 631898
rect 270804 596218 270986 596454
rect 271222 596218 271404 596454
rect 270804 596134 271404 596218
rect 270804 595898 270986 596134
rect 271222 595898 271404 596134
rect 262128 578454 262448 578476
rect 262128 578218 262170 578454
rect 262406 578218 262448 578454
rect 262128 578134 262448 578218
rect 262128 577898 262170 578134
rect 262406 577898 262448 578134
rect 262128 577876 262448 577898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 246768 560454 247088 560476
rect 246768 560218 246810 560454
rect 247046 560218 247088 560454
rect 246768 560134 247088 560218
rect 246768 559898 246810 560134
rect 247046 559898 247088 560134
rect 246768 559876 247088 559898
rect 270804 560454 271404 595898
rect 270804 560218 270986 560454
rect 271222 560218 271404 560454
rect 270804 560134 271404 560218
rect 270804 559898 270986 560134
rect 271222 559898 271404 560134
rect 262128 542454 262448 542476
rect 262128 542218 262170 542454
rect 262406 542218 262448 542454
rect 262128 542134 262448 542218
rect 262128 541898 262170 542134
rect 262406 541898 262448 542134
rect 262128 541876 262448 541898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 246768 524454 247088 524476
rect 246768 524218 246810 524454
rect 247046 524218 247088 524454
rect 246768 524134 247088 524218
rect 246768 523898 246810 524134
rect 247046 523898 247088 524134
rect 246768 523876 247088 523898
rect 270804 524454 271404 559898
rect 270804 524218 270986 524454
rect 271222 524218 271404 524454
rect 270804 524134 271404 524218
rect 270804 523898 270986 524134
rect 271222 523898 271404 524134
rect 262128 506454 262448 506476
rect 262128 506218 262170 506454
rect 262406 506218 262448 506454
rect 262128 506134 262448 506218
rect 262128 505898 262170 506134
rect 262406 505898 262448 506134
rect 262128 505876 262448 505898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 246768 488454 247088 488476
rect 246768 488218 246810 488454
rect 247046 488218 247088 488454
rect 246768 488134 247088 488218
rect 246768 487898 246810 488134
rect 247046 487898 247088 488134
rect 246768 487876 247088 487898
rect 270804 488454 271404 523898
rect 288804 704838 289404 705800
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 578454 289404 613898
rect 306804 705778 307404 705800
rect 306804 705542 306986 705778
rect 307222 705542 307404 705778
rect 306804 705458 307404 705542
rect 306804 705222 306986 705458
rect 307222 705222 307404 705458
rect 306804 668454 307404 705222
rect 324804 704838 325404 705800
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 310651 700228 310717 700229
rect 310651 700164 310652 700228
rect 310716 700164 310717 700228
rect 310651 700163 310717 700164
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 632454 307404 667898
rect 306804 632218 306986 632454
rect 307222 632218 307404 632454
rect 306804 632134 307404 632218
rect 306804 631898 306986 632134
rect 307222 631898 307404 632134
rect 306804 596454 307404 631898
rect 306804 596218 306986 596454
rect 307222 596218 307404 596454
rect 306804 596134 307404 596218
rect 306804 595898 306986 596134
rect 307222 595898 307404 596134
rect 306603 586532 306669 586533
rect 306603 586468 306604 586532
rect 306668 586468 306669 586532
rect 306603 586467 306669 586468
rect 289675 586260 289741 586261
rect 289675 586196 289676 586260
rect 289740 586196 289741 586260
rect 289675 586195 289741 586196
rect 289491 586124 289557 586125
rect 289491 586060 289492 586124
rect 289556 586060 289557 586124
rect 289491 586059 289557 586060
rect 288804 578218 288986 578454
rect 289222 578218 289404 578454
rect 288804 578134 289404 578218
rect 288804 577898 288986 578134
rect 289222 577898 289404 578134
rect 288804 542454 289404 577898
rect 288804 542218 288986 542454
rect 289222 542218 289404 542454
rect 288804 542134 289404 542218
rect 288804 541898 288986 542134
rect 289222 541898 289404 542134
rect 276427 510916 276493 510917
rect 276427 510852 276428 510916
rect 276492 510852 276493 510916
rect 276427 510851 276493 510852
rect 270804 488218 270986 488454
rect 271222 488218 271404 488454
rect 270804 488134 271404 488218
rect 270804 487898 270986 488134
rect 271222 487898 271404 488134
rect 262128 470454 262448 470476
rect 262128 470218 262170 470454
rect 262406 470218 262448 470454
rect 262128 470134 262448 470218
rect 262128 469898 262170 470134
rect 262406 469898 262448 470134
rect 262128 469876 262448 469898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 246768 452454 247088 452476
rect 246768 452218 246810 452454
rect 247046 452218 247088 452454
rect 246768 452134 247088 452218
rect 246768 451898 246810 452134
rect 247046 451898 247088 452134
rect 246768 451876 247088 451898
rect 270804 452454 271404 487898
rect 270804 452218 270986 452454
rect 271222 452218 271404 452454
rect 270804 452134 271404 452218
rect 270804 451898 270986 452134
rect 271222 451898 271404 452134
rect 262128 434454 262448 434476
rect 262128 434218 262170 434454
rect 262406 434218 262448 434454
rect 262128 434134 262448 434218
rect 262128 433898 262170 434134
rect 262406 433898 262448 434134
rect 262128 433876 262448 433898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 246768 416454 247088 416476
rect 246768 416218 246810 416454
rect 247046 416218 247088 416454
rect 246768 416134 247088 416218
rect 246768 415898 246810 416134
rect 247046 415898 247088 416134
rect 246768 415876 247088 415898
rect 270804 416454 271404 451898
rect 270804 416218 270986 416454
rect 271222 416218 271404 416454
rect 270804 416134 271404 416218
rect 270804 415898 270986 416134
rect 271222 415898 271404 416134
rect 262128 398454 262448 398476
rect 262128 398218 262170 398454
rect 262406 398218 262448 398454
rect 262128 398134 262448 398218
rect 262128 397898 262170 398134
rect 262406 397898 262448 398134
rect 262128 397876 262448 397898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 36804 362454 37404 382916
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 274600 37404 289898
rect 54804 380454 55404 382916
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 274600 55404 307898
rect 72804 362454 73404 382916
rect 72804 362218 72986 362454
rect 73222 362218 73404 362454
rect 72804 362134 73404 362218
rect 72804 361898 72986 362134
rect 73222 361898 73404 362134
rect 72804 326454 73404 361898
rect 72804 326218 72986 326454
rect 73222 326218 73404 326454
rect 72804 326134 73404 326218
rect 72804 325898 72986 326134
rect 73222 325898 73404 326134
rect 72804 290454 73404 325898
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 274600 73404 289898
rect 90804 380454 91404 382916
rect 90804 380218 90986 380454
rect 91222 380218 91404 380454
rect 90804 380134 91404 380218
rect 90804 379898 90986 380134
rect 91222 379898 91404 380134
rect 90804 344454 91404 379898
rect 90804 344218 90986 344454
rect 91222 344218 91404 344454
rect 90804 344134 91404 344218
rect 90804 343898 90986 344134
rect 91222 343898 91404 344134
rect 90804 308454 91404 343898
rect 90804 308218 90986 308454
rect 91222 308218 91404 308454
rect 90804 308134 91404 308218
rect 90804 307898 90986 308134
rect 91222 307898 91404 308134
rect 90804 274600 91404 307898
rect 108804 362454 109404 382916
rect 108804 362218 108986 362454
rect 109222 362218 109404 362454
rect 108804 362134 109404 362218
rect 108804 361898 108986 362134
rect 109222 361898 109404 362134
rect 108804 326454 109404 361898
rect 108804 326218 108986 326454
rect 109222 326218 109404 326454
rect 108804 326134 109404 326218
rect 108804 325898 108986 326134
rect 109222 325898 109404 326134
rect 108804 290454 109404 325898
rect 108804 290218 108986 290454
rect 109222 290218 109404 290454
rect 108804 290134 109404 290218
rect 108804 289898 108986 290134
rect 109222 289898 109404 290134
rect 108804 274600 109404 289898
rect 126804 380454 127404 382916
rect 126804 380218 126986 380454
rect 127222 380218 127404 380454
rect 126804 380134 127404 380218
rect 126804 379898 126986 380134
rect 127222 379898 127404 380134
rect 126804 344454 127404 379898
rect 126804 344218 126986 344454
rect 127222 344218 127404 344454
rect 126804 344134 127404 344218
rect 126804 343898 126986 344134
rect 127222 343898 127404 344134
rect 126804 308454 127404 343898
rect 126804 308218 126986 308454
rect 127222 308218 127404 308454
rect 126804 308134 127404 308218
rect 126804 307898 126986 308134
rect 127222 307898 127404 308134
rect 126804 274600 127404 307898
rect 144804 362454 145404 382916
rect 144804 362218 144986 362454
rect 145222 362218 145404 362454
rect 144804 362134 145404 362218
rect 144804 361898 144986 362134
rect 145222 361898 145404 362134
rect 144804 326454 145404 361898
rect 144804 326218 144986 326454
rect 145222 326218 145404 326454
rect 144804 326134 145404 326218
rect 144804 325898 144986 326134
rect 145222 325898 145404 326134
rect 144804 290454 145404 325898
rect 144804 290218 144986 290454
rect 145222 290218 145404 290454
rect 144804 290134 145404 290218
rect 144804 289898 144986 290134
rect 145222 289898 145404 290134
rect 144804 274600 145404 289898
rect 162804 380454 163404 382916
rect 162804 380218 162986 380454
rect 163222 380218 163404 380454
rect 162804 380134 163404 380218
rect 162804 379898 162986 380134
rect 163222 379898 163404 380134
rect 162804 344454 163404 379898
rect 162804 344218 162986 344454
rect 163222 344218 163404 344454
rect 162804 344134 163404 344218
rect 162804 343898 162986 344134
rect 163222 343898 163404 344134
rect 162804 308454 163404 343898
rect 162804 308218 162986 308454
rect 163222 308218 163404 308454
rect 162804 308134 163404 308218
rect 162804 307898 162986 308134
rect 163222 307898 163404 308134
rect 162804 274600 163404 307898
rect 180804 362454 181404 382916
rect 180804 362218 180986 362454
rect 181222 362218 181404 362454
rect 180804 362134 181404 362218
rect 180804 361898 180986 362134
rect 181222 361898 181404 362134
rect 180804 326454 181404 361898
rect 180804 326218 180986 326454
rect 181222 326218 181404 326454
rect 180804 326134 181404 326218
rect 180804 325898 180986 326134
rect 181222 325898 181404 326134
rect 180804 290454 181404 325898
rect 180804 290218 180986 290454
rect 181222 290218 181404 290454
rect 180804 290134 181404 290218
rect 180804 289898 180986 290134
rect 181222 289898 181404 290134
rect 180804 274600 181404 289898
rect 198804 380454 199404 382916
rect 198804 380218 198986 380454
rect 199222 380218 199404 380454
rect 198804 380134 199404 380218
rect 198804 379898 198986 380134
rect 199222 379898 199404 380134
rect 198804 344454 199404 379898
rect 198804 344218 198986 344454
rect 199222 344218 199404 344454
rect 198804 344134 199404 344218
rect 198804 343898 198986 344134
rect 199222 343898 199404 344134
rect 198804 308454 199404 343898
rect 198804 308218 198986 308454
rect 199222 308218 199404 308454
rect 198804 308134 199404 308218
rect 198804 307898 198986 308134
rect 199222 307898 199404 308134
rect 198804 274600 199404 307898
rect 216804 362454 217404 382916
rect 216804 362218 216986 362454
rect 217222 362218 217404 362454
rect 216804 362134 217404 362218
rect 216804 361898 216986 362134
rect 217222 361898 217404 362134
rect 216804 326454 217404 361898
rect 216804 326218 216986 326454
rect 217222 326218 217404 326454
rect 216804 326134 217404 326218
rect 216804 325898 216986 326134
rect 217222 325898 217404 326134
rect 216804 290454 217404 325898
rect 216804 290218 216986 290454
rect 217222 290218 217404 290454
rect 216804 290134 217404 290218
rect 216804 289898 216986 290134
rect 217222 289898 217404 290134
rect 216804 274600 217404 289898
rect 234804 380454 235404 382916
rect 234804 380218 234986 380454
rect 235222 380218 235404 380454
rect 234804 380134 235404 380218
rect 234804 379898 234986 380134
rect 235222 379898 235404 380134
rect 234804 344454 235404 379898
rect 234804 344218 234986 344454
rect 235222 344218 235404 344454
rect 234804 344134 235404 344218
rect 234804 343898 234986 344134
rect 235222 343898 235404 344134
rect 234804 308454 235404 343898
rect 234804 308218 234986 308454
rect 235222 308218 235404 308454
rect 234804 308134 235404 308218
rect 234804 307898 234986 308134
rect 235222 307898 235404 308134
rect 234804 274600 235404 307898
rect 252804 362454 253404 382916
rect 252804 362218 252986 362454
rect 253222 362218 253404 362454
rect 252804 362134 253404 362218
rect 252804 361898 252986 362134
rect 253222 361898 253404 362134
rect 252804 326454 253404 361898
rect 270804 380454 271404 415898
rect 275139 382260 275205 382261
rect 275139 382196 275140 382260
rect 275204 382196 275205 382260
rect 275139 382195 275205 382196
rect 274955 381988 275021 381989
rect 274955 381924 274956 381988
rect 275020 381924 275021 381988
rect 274955 381923 275021 381924
rect 270804 380218 270986 380454
rect 271222 380218 271404 380454
rect 270804 380134 271404 380218
rect 270804 379898 270986 380134
rect 271222 379898 271404 380134
rect 270804 356560 271404 379898
rect 252804 326218 252986 326454
rect 253222 326218 253404 326454
rect 252804 326134 253404 326218
rect 252804 325898 252986 326134
rect 253222 325898 253404 326134
rect 252804 290454 253404 325898
rect 252804 290218 252986 290454
rect 253222 290218 253404 290454
rect 252804 290134 253404 290218
rect 252804 289898 252986 290134
rect 253222 289898 253404 290134
rect 252804 274600 253404 289898
rect 270804 308454 271404 314560
rect 274958 313173 275018 381923
rect 275142 313309 275202 382195
rect 275875 354924 275941 354925
rect 275875 354860 275876 354924
rect 275940 354860 275941 354924
rect 275875 354859 275941 354860
rect 275139 313308 275205 313309
rect 275139 313244 275140 313308
rect 275204 313244 275205 313308
rect 275139 313243 275205 313244
rect 274955 313172 275021 313173
rect 274955 313108 274956 313172
rect 275020 313108 275021 313172
rect 274955 313107 275021 313108
rect 270804 308218 270986 308454
rect 271222 308218 271404 308454
rect 270804 308134 271404 308218
rect 270804 307898 270986 308134
rect 271222 307898 271404 308134
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 270804 272454 271404 307898
rect 275878 273733 275938 354859
rect 276430 315621 276490 510851
rect 288804 506454 289404 541898
rect 288804 506218 288986 506454
rect 289222 506218 289404 506454
rect 288804 506134 289404 506218
rect 288804 505898 288986 506134
rect 289222 505898 289404 506134
rect 288804 470454 289404 505898
rect 288804 470218 288986 470454
rect 289222 470218 289404 470454
rect 288804 470134 289404 470218
rect 288804 469898 288986 470134
rect 289222 469898 289404 470134
rect 288804 434454 289404 469898
rect 288804 434218 288986 434454
rect 289222 434218 289404 434454
rect 288804 434134 289404 434218
rect 288804 433898 288986 434134
rect 289222 433898 289404 434134
rect 288804 398454 289404 433898
rect 288804 398218 288986 398454
rect 289222 398218 289404 398454
rect 288804 398134 289404 398218
rect 288804 397898 288986 398134
rect 289222 397898 289404 398134
rect 288804 362454 289404 397898
rect 288804 362218 288986 362454
rect 289222 362218 289404 362454
rect 288804 362134 289404 362218
rect 288804 361898 288986 362134
rect 289222 361898 289404 362134
rect 276611 359276 276677 359277
rect 276611 359212 276612 359276
rect 276676 359212 276677 359276
rect 276611 359211 276677 359212
rect 276427 315620 276493 315621
rect 276427 315556 276428 315620
rect 276492 315556 276493 315620
rect 276427 315555 276493 315556
rect 275875 273732 275941 273733
rect 275875 273668 275876 273732
rect 275940 273668 275941 273732
rect 275875 273667 275941 273668
rect 270804 272218 270986 272454
rect 271222 272218 271404 272454
rect 270804 272134 271404 272218
rect 270804 271898 270986 272134
rect 271222 271898 271404 272134
rect 262128 254454 262448 254476
rect 262128 254218 262170 254454
rect 262406 254218 262448 254454
rect 262128 254134 262448 254218
rect 262128 253898 262170 254134
rect 262406 253898 262448 254134
rect 262128 253876 262448 253898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 246768 236454 247088 236476
rect 246768 236218 246810 236454
rect 247046 236218 247088 236454
rect 246768 236134 247088 236218
rect 246768 235898 246810 236134
rect 247046 235898 247088 236134
rect 246768 235876 247088 235898
rect 270804 236454 271404 271898
rect 270804 236218 270986 236454
rect 271222 236218 271404 236454
rect 270804 236134 271404 236218
rect 270804 235898 270986 236134
rect 271222 235898 271404 236134
rect 262128 218454 262448 218476
rect 262128 218218 262170 218454
rect 262406 218218 262448 218454
rect 262128 218134 262448 218218
rect 262128 217898 262170 218134
rect 262406 217898 262448 218134
rect 262128 217876 262448 217898
rect 270171 216340 270237 216341
rect 270171 216276 270172 216340
rect 270236 216276 270237 216340
rect 270171 216275 270237 216276
rect 270174 206141 270234 216275
rect 270171 206140 270237 206141
rect 270171 206076 270172 206140
rect 270236 206076 270237 206140
rect 270171 206075 270237 206076
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 246768 200454 247088 200476
rect 246768 200218 246810 200454
rect 247046 200218 247088 200454
rect 246768 200134 247088 200218
rect 246768 199898 246810 200134
rect 247046 199898 247088 200134
rect 246768 199876 247088 199898
rect 270804 200454 271404 235898
rect 270804 200218 270986 200454
rect 271222 200218 271404 200454
rect 270804 200134 271404 200218
rect 270804 199898 270986 200134
rect 271222 199898 271404 200134
rect 262128 182454 262448 182476
rect 262128 182218 262170 182454
rect 262406 182218 262448 182454
rect 262128 182134 262448 182218
rect 262128 181898 262170 182134
rect 262406 181898 262448 182134
rect 262128 181876 262448 181898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 246768 164454 247088 164476
rect 246768 164218 246810 164454
rect 247046 164218 247088 164454
rect 246768 164134 247088 164218
rect 246768 163898 246810 164134
rect 247046 163898 247088 164134
rect 246768 163876 247088 163898
rect 270804 164454 271404 199898
rect 270804 164218 270986 164454
rect 271222 164218 271404 164454
rect 270804 164134 271404 164218
rect 270804 163898 270986 164134
rect 271222 163898 271404 164134
rect 262128 146454 262448 146476
rect 262128 146218 262170 146454
rect 262406 146218 262448 146454
rect 262128 146134 262448 146218
rect 262128 145898 262170 146134
rect 262406 145898 262448 146134
rect 262128 145876 262448 145898
rect 270171 134060 270237 134061
rect 270171 133996 270172 134060
rect 270236 133996 270237 134060
rect 270171 133995 270237 133996
rect 270174 132565 270234 133995
rect 270171 132564 270237 132565
rect 270171 132500 270172 132564
rect 270236 132500 270237 132564
rect 270171 132499 270237 132500
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 246768 128454 247088 128476
rect 246768 128218 246810 128454
rect 247046 128218 247088 128454
rect 246768 128134 247088 128218
rect 246768 127898 246810 128134
rect 247046 127898 247088 128134
rect 246768 127876 247088 127898
rect 270804 128454 271404 163898
rect 270804 128218 270986 128454
rect 271222 128218 271404 128454
rect 270804 128134 271404 128218
rect 270804 127898 270986 128134
rect 271222 127898 271404 128134
rect 262128 110454 262448 110476
rect 262128 110218 262170 110454
rect 262406 110218 262448 110454
rect 262128 110134 262448 110218
rect 262128 109898 262170 110134
rect 262406 109898 262448 110134
rect 262128 109876 262448 109898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 246768 92454 247088 92476
rect 246768 92218 246810 92454
rect 247046 92218 247088 92454
rect 246768 92134 247088 92218
rect 246768 91898 246810 92134
rect 247046 91898 247088 92134
rect 246768 91876 247088 91898
rect 270804 92454 271404 127898
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1286 19404 19898
rect 18804 -1522 18986 -1286
rect 19222 -1522 19404 -1286
rect 18804 -1606 19404 -1522
rect 18804 -1842 18986 -1606
rect 19222 -1842 19404 -1606
rect 18804 -1864 19404 -1842
rect 36804 38454 37404 72600
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1864 37404 -902
rect 54804 56454 55404 72600
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1286 55404 19898
rect 54804 -1522 54986 -1286
rect 55222 -1522 55404 -1286
rect 54804 -1606 55404 -1522
rect 54804 -1842 54986 -1606
rect 55222 -1842 55404 -1606
rect 54804 -1864 55404 -1842
rect 72804 38454 73404 72600
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1864 73404 -902
rect 90804 56454 91404 72600
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1286 91404 19898
rect 90804 -1522 90986 -1286
rect 91222 -1522 91404 -1286
rect 90804 -1606 91404 -1522
rect 90804 -1842 90986 -1606
rect 91222 -1842 91404 -1606
rect 90804 -1864 91404 -1842
rect 108804 38454 109404 72600
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1864 109404 -902
rect 126804 56454 127404 72600
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1286 127404 19898
rect 126804 -1522 126986 -1286
rect 127222 -1522 127404 -1286
rect 126804 -1606 127404 -1522
rect 126804 -1842 126986 -1606
rect 127222 -1842 127404 -1606
rect 126804 -1864 127404 -1842
rect 144804 38454 145404 72600
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1864 145404 -902
rect 162804 56454 163404 72600
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1286 163404 19898
rect 162804 -1522 162986 -1286
rect 163222 -1522 163404 -1286
rect 162804 -1606 163404 -1522
rect 162804 -1842 162986 -1606
rect 163222 -1842 163404 -1606
rect 162804 -1864 163404 -1842
rect 180804 38454 181404 72600
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1864 181404 -902
rect 198804 56454 199404 72600
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1286 199404 19898
rect 198804 -1522 198986 -1286
rect 199222 -1522 199404 -1286
rect 198804 -1606 199404 -1522
rect 198804 -1842 198986 -1606
rect 199222 -1842 199404 -1606
rect 198804 -1864 199404 -1842
rect 216804 38454 217404 72600
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1864 217404 -902
rect 234804 56454 235404 72600
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 234804 20454 235404 55898
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1286 235404 19898
rect 234804 -1522 234986 -1286
rect 235222 -1522 235404 -1286
rect 234804 -1606 235404 -1522
rect 234804 -1842 234986 -1606
rect 235222 -1842 235404 -1606
rect 234804 -1864 235404 -1842
rect 252804 38454 253404 72600
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1864 253404 -902
rect 270804 56454 271404 91898
rect 276614 72045 276674 359211
rect 288804 356560 289404 361898
rect 287835 354924 287901 354925
rect 287835 354860 287836 354924
rect 287900 354860 287901 354924
rect 287835 354859 287901 354860
rect 287838 133925 287898 354859
rect 288804 290454 289404 314560
rect 289494 313309 289554 586059
rect 289678 313445 289738 586195
rect 298691 586124 298757 586125
rect 298691 586060 298692 586124
rect 298756 586060 298757 586124
rect 298691 586059 298757 586060
rect 297219 382124 297285 382125
rect 297219 382060 297220 382124
rect 297284 382060 297285 382124
rect 297219 382059 297285 382060
rect 289859 354924 289925 354925
rect 289859 354860 289860 354924
rect 289924 354860 289925 354924
rect 289859 354859 289925 354860
rect 291331 354924 291397 354925
rect 291331 354860 291332 354924
rect 291396 354860 291397 354924
rect 291331 354859 291397 354860
rect 293539 354924 293605 354925
rect 293539 354860 293540 354924
rect 293604 354860 293605 354924
rect 293539 354859 293605 354860
rect 289675 313444 289741 313445
rect 289675 313380 289676 313444
rect 289740 313380 289741 313444
rect 289675 313379 289741 313380
rect 289491 313308 289557 313309
rect 289491 313244 289492 313308
rect 289556 313244 289557 313308
rect 289491 313243 289557 313244
rect 288804 290218 288986 290454
rect 289222 290218 289404 290454
rect 288804 290134 289404 290218
rect 288804 289898 288986 290134
rect 289222 289898 289404 290134
rect 288804 254454 289404 289898
rect 289862 276725 289922 354859
rect 289859 276724 289925 276725
rect 289859 276660 289860 276724
rect 289924 276660 289925 276724
rect 289859 276659 289925 276660
rect 291334 276045 291394 354859
rect 292112 344454 292432 344476
rect 292112 344218 292154 344454
rect 292390 344218 292432 344454
rect 292112 344134 292432 344218
rect 292112 343898 292154 344134
rect 292390 343898 292432 344134
rect 292112 343876 292432 343898
rect 293542 276725 293602 354859
rect 297222 316301 297282 382059
rect 298694 316301 298754 586059
rect 304579 385660 304645 385661
rect 304579 385596 304580 385660
rect 304644 385596 304645 385660
rect 304579 385595 304645 385596
rect 300899 354924 300965 354925
rect 300899 354860 300900 354924
rect 300964 354860 300965 354924
rect 300899 354859 300965 354860
rect 297219 316300 297285 316301
rect 297219 316236 297220 316300
rect 297284 316236 297285 316300
rect 297219 316235 297285 316236
rect 298691 316300 298757 316301
rect 298691 316236 298692 316300
rect 298756 316236 298757 316300
rect 298691 316235 298757 316236
rect 293539 276724 293605 276725
rect 293539 276660 293540 276724
rect 293604 276660 293605 276724
rect 293539 276659 293605 276660
rect 291331 276044 291397 276045
rect 291331 275980 291332 276044
rect 291396 275980 291397 276044
rect 291331 275979 291397 275980
rect 288804 254218 288986 254454
rect 289222 254218 289404 254454
rect 288804 254134 289404 254218
rect 288804 253898 288986 254134
rect 289222 253898 289404 254134
rect 288804 218454 289404 253898
rect 288804 218218 288986 218454
rect 289222 218218 289404 218454
rect 288804 218134 289404 218218
rect 288804 217898 288986 218134
rect 289222 217898 289404 218134
rect 288804 182454 289404 217898
rect 288804 182218 288986 182454
rect 289222 182218 289404 182454
rect 288804 182134 289404 182218
rect 288804 181898 288986 182134
rect 289222 181898 289404 182134
rect 288804 146454 289404 181898
rect 288804 146218 288986 146454
rect 289222 146218 289404 146454
rect 288804 146134 289404 146218
rect 288804 145898 288986 146134
rect 289222 145898 289404 146134
rect 287835 133924 287901 133925
rect 287835 133860 287836 133924
rect 287900 133860 287901 133924
rect 287835 133859 287901 133860
rect 288804 110454 289404 145898
rect 288804 110218 288986 110454
rect 289222 110218 289404 110454
rect 288804 110134 289404 110218
rect 288804 109898 288986 110134
rect 289222 109898 289404 110134
rect 288804 74454 289404 109898
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 276611 72044 276677 72045
rect 276611 71980 276612 72044
rect 276676 71980 276677 72044
rect 276611 71979 276677 71980
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1286 271404 19898
rect 270804 -1522 270986 -1286
rect 271222 -1522 271404 -1286
rect 270804 -1606 271404 -1522
rect 270804 -1842 270986 -1606
rect 271222 -1842 271404 -1606
rect 270804 -1864 271404 -1842
rect 288804 38454 289404 73898
rect 300902 72045 300962 354859
rect 304582 315485 304642 385595
rect 306419 354924 306485 354925
rect 306419 354860 306420 354924
rect 306484 354860 306485 354924
rect 306419 354859 306485 354860
rect 304579 315484 304645 315485
rect 304579 315420 304580 315484
rect 304644 315420 304645 315484
rect 304579 315419 304645 315420
rect 306422 272237 306482 354859
rect 306606 315621 306666 586467
rect 306804 560454 307404 595898
rect 306804 560218 306986 560454
rect 307222 560218 307404 560454
rect 306804 560134 307404 560218
rect 306804 559898 306986 560134
rect 307222 559898 307404 560134
rect 306804 524454 307404 559898
rect 306804 524218 306986 524454
rect 307222 524218 307404 524454
rect 306804 524134 307404 524218
rect 306804 523898 306986 524134
rect 307222 523898 307404 524134
rect 306804 488454 307404 523898
rect 306804 488218 306986 488454
rect 307222 488218 307404 488454
rect 306804 488134 307404 488218
rect 306804 487898 306986 488134
rect 307222 487898 307404 488134
rect 306804 452454 307404 487898
rect 306804 452218 306986 452454
rect 307222 452218 307404 452454
rect 306804 452134 307404 452218
rect 306804 451898 306986 452134
rect 307222 451898 307404 452134
rect 306804 416454 307404 451898
rect 306804 416218 306986 416454
rect 307222 416218 307404 416454
rect 306804 416134 307404 416218
rect 306804 415898 306986 416134
rect 307222 415898 307404 416134
rect 306804 380454 307404 415898
rect 306804 380218 306986 380454
rect 307222 380218 307404 380454
rect 306804 380134 307404 380218
rect 306804 379898 306986 380134
rect 307222 379898 307404 380134
rect 306804 356560 307404 379898
rect 307472 326454 307792 326476
rect 307472 326218 307514 326454
rect 307750 326218 307792 326454
rect 307472 326134 307792 326218
rect 307472 325898 307514 326134
rect 307750 325898 307792 326134
rect 307472 325876 307792 325898
rect 310654 318610 310714 700163
rect 311019 700092 311085 700093
rect 311019 700028 311020 700092
rect 311084 700028 311085 700092
rect 311019 700027 311085 700028
rect 310835 699956 310901 699957
rect 310835 699892 310836 699956
rect 310900 699892 310901 699956
rect 310835 699891 310901 699892
rect 310838 322010 310898 699891
rect 311022 324730 311082 700027
rect 311939 699956 312005 699957
rect 311939 699892 311940 699956
rect 312004 699892 312005 699956
rect 311939 699891 312005 699892
rect 311203 585988 311269 585989
rect 311203 585924 311204 585988
rect 311268 585924 311269 585988
rect 311203 585923 311269 585924
rect 311206 343090 311266 585923
rect 311571 343092 311637 343093
rect 311571 343090 311572 343092
rect 311206 343030 311572 343090
rect 311571 343028 311572 343030
rect 311636 343028 311637 343092
rect 311571 343027 311637 343028
rect 311571 324732 311637 324733
rect 311571 324730 311572 324732
rect 311022 324670 311572 324730
rect 311571 324668 311572 324670
rect 311636 324668 311637 324732
rect 311571 324667 311637 324668
rect 311571 322012 311637 322013
rect 311571 322010 311572 322012
rect 310838 321950 311572 322010
rect 311571 321948 311572 321950
rect 311636 321948 311637 322012
rect 311571 321947 311637 321948
rect 311571 318612 311637 318613
rect 311571 318610 311572 318612
rect 310654 318550 311572 318610
rect 311571 318548 311572 318550
rect 311636 318548 311637 318612
rect 311571 318547 311637 318548
rect 311942 316301 312002 699891
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 650454 325404 685898
rect 324804 650218 324986 650454
rect 325222 650218 325404 650454
rect 324804 650134 325404 650218
rect 324804 649898 324986 650134
rect 325222 649898 325404 650134
rect 324804 614454 325404 649898
rect 324804 614218 324986 614454
rect 325222 614218 325404 614454
rect 324804 614134 325404 614218
rect 324804 613898 324986 614134
rect 325222 613898 325404 614134
rect 324804 584916 325404 613898
rect 342804 705778 343404 705800
rect 342804 705542 342986 705778
rect 343222 705542 343404 705778
rect 342804 705458 343404 705542
rect 342804 705222 342986 705458
rect 343222 705222 343404 705458
rect 342804 668454 343404 705222
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 632454 343404 667898
rect 342804 632218 342986 632454
rect 343222 632218 343404 632454
rect 342804 632134 343404 632218
rect 342804 631898 342986 632134
rect 343222 631898 343404 632134
rect 342804 596454 343404 631898
rect 342804 596218 342986 596454
rect 343222 596218 343404 596454
rect 342804 596134 343404 596218
rect 342804 595898 342986 596134
rect 343222 595898 343404 596134
rect 342804 584916 343404 595898
rect 360804 704838 361404 705800
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 650454 361404 685898
rect 360804 650218 360986 650454
rect 361222 650218 361404 650454
rect 360804 650134 361404 650218
rect 360804 649898 360986 650134
rect 361222 649898 361404 650134
rect 360804 614454 361404 649898
rect 360804 614218 360986 614454
rect 361222 614218 361404 614454
rect 360804 614134 361404 614218
rect 360804 613898 360986 614134
rect 361222 613898 361404 614134
rect 360804 584916 361404 613898
rect 378804 705778 379404 705800
rect 378804 705542 378986 705778
rect 379222 705542 379404 705778
rect 378804 705458 379404 705542
rect 378804 705222 378986 705458
rect 379222 705222 379404 705458
rect 378804 668454 379404 705222
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 632454 379404 667898
rect 378804 632218 378986 632454
rect 379222 632218 379404 632454
rect 378804 632134 379404 632218
rect 378804 631898 378986 632134
rect 379222 631898 379404 632134
rect 378804 596454 379404 631898
rect 378804 596218 378986 596454
rect 379222 596218 379404 596454
rect 378804 596134 379404 596218
rect 378804 595898 378986 596134
rect 379222 595898 379404 596134
rect 378804 584916 379404 595898
rect 396804 704838 397404 705800
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 396804 614454 397404 649898
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 396804 584916 397404 613898
rect 414804 705778 415404 705800
rect 414804 705542 414986 705778
rect 415222 705542 415404 705778
rect 414804 705458 415404 705542
rect 414804 705222 414986 705458
rect 415222 705222 415404 705458
rect 414804 668454 415404 705222
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 632454 415404 667898
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 596454 415404 631898
rect 414804 596218 414986 596454
rect 415222 596218 415404 596454
rect 414804 596134 415404 596218
rect 414804 595898 414986 596134
rect 415222 595898 415404 596134
rect 414804 584916 415404 595898
rect 432804 704838 433404 705800
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 614454 433404 649898
rect 432804 614218 432986 614454
rect 433222 614218 433404 614454
rect 432804 614134 433404 614218
rect 432804 613898 432986 614134
rect 433222 613898 433404 614134
rect 432804 584916 433404 613898
rect 450804 705778 451404 705800
rect 450804 705542 450986 705778
rect 451222 705542 451404 705778
rect 450804 705458 451404 705542
rect 450804 705222 450986 705458
rect 451222 705222 451404 705458
rect 450804 668454 451404 705222
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 632454 451404 667898
rect 450804 632218 450986 632454
rect 451222 632218 451404 632454
rect 450804 632134 451404 632218
rect 450804 631898 450986 632134
rect 451222 631898 451404 632134
rect 450804 596454 451404 631898
rect 450804 596218 450986 596454
rect 451222 596218 451404 596454
rect 450804 596134 451404 596218
rect 450804 595898 450986 596134
rect 451222 595898 451404 596134
rect 450804 584916 451404 595898
rect 468804 704838 469404 705800
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 650454 469404 685898
rect 468804 650218 468986 650454
rect 469222 650218 469404 650454
rect 468804 650134 469404 650218
rect 468804 649898 468986 650134
rect 469222 649898 469404 650134
rect 468804 614454 469404 649898
rect 468804 614218 468986 614454
rect 469222 614218 469404 614454
rect 468804 614134 469404 614218
rect 468804 613898 468986 614134
rect 469222 613898 469404 614134
rect 468804 584916 469404 613898
rect 486804 705778 487404 705800
rect 486804 705542 486986 705778
rect 487222 705542 487404 705778
rect 486804 705458 487404 705542
rect 486804 705222 486986 705458
rect 487222 705222 487404 705458
rect 486804 668454 487404 705222
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 632454 487404 667898
rect 486804 632218 486986 632454
rect 487222 632218 487404 632454
rect 486804 632134 487404 632218
rect 486804 631898 486986 632134
rect 487222 631898 487404 632134
rect 486804 596454 487404 631898
rect 486804 596218 486986 596454
rect 487222 596218 487404 596454
rect 486804 596134 487404 596218
rect 486804 595898 486986 596134
rect 487222 595898 487404 596134
rect 486804 584916 487404 595898
rect 504804 704838 505404 705800
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 650454 505404 685898
rect 504804 650218 504986 650454
rect 505222 650218 505404 650454
rect 504804 650134 505404 650218
rect 504804 649898 504986 650134
rect 505222 649898 505404 650134
rect 504804 614454 505404 649898
rect 504804 614218 504986 614454
rect 505222 614218 505404 614454
rect 504804 614134 505404 614218
rect 504804 613898 504986 614134
rect 505222 613898 505404 614134
rect 504804 584916 505404 613898
rect 522804 705778 523404 705800
rect 522804 705542 522986 705778
rect 523222 705542 523404 705778
rect 522804 705458 523404 705542
rect 522804 705222 522986 705458
rect 523222 705222 523404 705458
rect 522804 668454 523404 705222
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522804 584916 523404 595898
rect 540804 704838 541404 705800
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 584916 541404 613898
rect 558804 705778 559404 705800
rect 558804 705542 558986 705778
rect 559222 705542 559404 705778
rect 558804 705458 559404 705542
rect 558804 705222 558986 705458
rect 559222 705222 559404 705458
rect 558804 668454 559404 705222
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 584916 559404 595898
rect 576804 704838 577404 705800
rect 586260 705778 586860 705800
rect 586260 705542 586442 705778
rect 586678 705542 586860 705778
rect 586260 705458 586860 705542
rect 586260 705222 586442 705458
rect 586678 705222 586860 705458
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 554256 578454 554576 578476
rect 554256 578218 554298 578454
rect 554534 578218 554576 578454
rect 554256 578134 554576 578218
rect 554256 577898 554298 578134
rect 554534 577898 554576 578134
rect 554256 577876 554576 577898
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 314147 565180 314213 565181
rect 314147 565116 314148 565180
rect 314212 565116 314213 565180
rect 314147 565115 314213 565116
rect 314150 559333 314210 565115
rect 538896 560454 539216 560476
rect 538896 560218 538938 560454
rect 539174 560218 539216 560454
rect 538896 560134 539216 560218
rect 538896 559898 538938 560134
rect 539174 559898 539216 560134
rect 538896 559876 539216 559898
rect 314147 559332 314213 559333
rect 314147 559268 314148 559332
rect 314212 559268 314213 559332
rect 314147 559267 314213 559268
rect 554256 542454 554576 542476
rect 554256 542218 554298 542454
rect 554534 542218 554576 542454
rect 554256 542134 554576 542218
rect 554256 541898 554298 542134
rect 554534 541898 554576 542134
rect 554256 541876 554576 541898
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 538896 524454 539216 524476
rect 538896 524218 538938 524454
rect 539174 524218 539216 524454
rect 538896 524134 539216 524218
rect 538896 523898 538938 524134
rect 539174 523898 539216 524134
rect 538896 523876 539216 523898
rect 554256 506454 554576 506476
rect 554256 506218 554298 506454
rect 554534 506218 554576 506454
rect 554256 506134 554576 506218
rect 554256 505898 554298 506134
rect 554534 505898 554576 506134
rect 554256 505876 554576 505898
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 538896 488454 539216 488476
rect 538896 488218 538938 488454
rect 539174 488218 539216 488454
rect 538896 488134 539216 488218
rect 538896 487898 538938 488134
rect 539174 487898 539216 488134
rect 538896 487876 539216 487898
rect 554256 470454 554576 470476
rect 554256 470218 554298 470454
rect 554534 470218 554576 470454
rect 554256 470134 554576 470218
rect 554256 469898 554298 470134
rect 554534 469898 554576 470134
rect 554256 469876 554576 469898
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 538896 452454 539216 452476
rect 538896 452218 538938 452454
rect 539174 452218 539216 452454
rect 538896 452134 539216 452218
rect 538896 451898 538938 452134
rect 539174 451898 539216 452134
rect 538896 451876 539216 451898
rect 554256 434454 554576 434476
rect 554256 434218 554298 434454
rect 554534 434218 554576 434454
rect 554256 434134 554576 434218
rect 554256 433898 554298 434134
rect 554534 433898 554576 434134
rect 554256 433876 554576 433898
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 538896 416454 539216 416476
rect 538896 416218 538938 416454
rect 539174 416218 539216 416454
rect 538896 416134 539216 416218
rect 538896 415898 538938 416134
rect 539174 415898 539216 416134
rect 538896 415876 539216 415898
rect 554256 398454 554576 398476
rect 554256 398218 554298 398454
rect 554534 398218 554576 398454
rect 554256 398134 554576 398218
rect 554256 397898 554298 398134
rect 554534 397898 554576 398134
rect 554256 397876 554576 397898
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 324804 362454 325404 382916
rect 324804 362218 324986 362454
rect 325222 362218 325404 362454
rect 324804 362134 325404 362218
rect 324804 361898 324986 362134
rect 325222 361898 325404 362134
rect 324804 326454 325404 361898
rect 324804 326218 324986 326454
rect 325222 326218 325404 326454
rect 324804 326134 325404 326218
rect 324804 325898 324986 326134
rect 325222 325898 325404 326134
rect 311939 316300 312005 316301
rect 311939 316236 311940 316300
rect 312004 316236 312005 316300
rect 311939 316235 312005 316236
rect 306603 315620 306669 315621
rect 306603 315556 306604 315620
rect 306668 315556 306669 315620
rect 306603 315555 306669 315556
rect 306804 308454 307404 314560
rect 306804 308218 306986 308454
rect 307222 308218 307404 308454
rect 306804 308134 307404 308218
rect 306804 307898 306986 308134
rect 307222 307898 307404 308134
rect 306804 272454 307404 307898
rect 324804 290454 325404 325898
rect 324804 290218 324986 290454
rect 325222 290218 325404 290454
rect 324804 290134 325404 290218
rect 324804 289898 324986 290134
rect 325222 289898 325404 290134
rect 324804 274600 325404 289898
rect 342804 380454 343404 382916
rect 342804 380218 342986 380454
rect 343222 380218 343404 380454
rect 342804 380134 343404 380218
rect 342804 379898 342986 380134
rect 343222 379898 343404 380134
rect 342804 344454 343404 379898
rect 342804 344218 342986 344454
rect 343222 344218 343404 344454
rect 342804 344134 343404 344218
rect 342804 343898 342986 344134
rect 343222 343898 343404 344134
rect 342804 308454 343404 343898
rect 342804 308218 342986 308454
rect 343222 308218 343404 308454
rect 342804 308134 343404 308218
rect 342804 307898 342986 308134
rect 343222 307898 343404 308134
rect 342804 274600 343404 307898
rect 360804 362454 361404 382916
rect 360804 362218 360986 362454
rect 361222 362218 361404 362454
rect 360804 362134 361404 362218
rect 360804 361898 360986 362134
rect 361222 361898 361404 362134
rect 360804 326454 361404 361898
rect 360804 326218 360986 326454
rect 361222 326218 361404 326454
rect 360804 326134 361404 326218
rect 360804 325898 360986 326134
rect 361222 325898 361404 326134
rect 360804 290454 361404 325898
rect 360804 290218 360986 290454
rect 361222 290218 361404 290454
rect 360804 290134 361404 290218
rect 360804 289898 360986 290134
rect 361222 289898 361404 290134
rect 360804 274600 361404 289898
rect 378804 380454 379404 382916
rect 378804 380218 378986 380454
rect 379222 380218 379404 380454
rect 378804 380134 379404 380218
rect 378804 379898 378986 380134
rect 379222 379898 379404 380134
rect 378804 344454 379404 379898
rect 378804 344218 378986 344454
rect 379222 344218 379404 344454
rect 378804 344134 379404 344218
rect 378804 343898 378986 344134
rect 379222 343898 379404 344134
rect 378804 308454 379404 343898
rect 378804 308218 378986 308454
rect 379222 308218 379404 308454
rect 378804 308134 379404 308218
rect 378804 307898 378986 308134
rect 379222 307898 379404 308134
rect 378804 274600 379404 307898
rect 396804 362454 397404 382916
rect 396804 362218 396986 362454
rect 397222 362218 397404 362454
rect 396804 362134 397404 362218
rect 396804 361898 396986 362134
rect 397222 361898 397404 362134
rect 396804 326454 397404 361898
rect 396804 326218 396986 326454
rect 397222 326218 397404 326454
rect 396804 326134 397404 326218
rect 396804 325898 396986 326134
rect 397222 325898 397404 326134
rect 396804 290454 397404 325898
rect 396804 290218 396986 290454
rect 397222 290218 397404 290454
rect 396804 290134 397404 290218
rect 396804 289898 396986 290134
rect 397222 289898 397404 290134
rect 396804 274600 397404 289898
rect 414804 380454 415404 382916
rect 414804 380218 414986 380454
rect 415222 380218 415404 380454
rect 414804 380134 415404 380218
rect 414804 379898 414986 380134
rect 415222 379898 415404 380134
rect 414804 344454 415404 379898
rect 414804 344218 414986 344454
rect 415222 344218 415404 344454
rect 414804 344134 415404 344218
rect 414804 343898 414986 344134
rect 415222 343898 415404 344134
rect 414804 308454 415404 343898
rect 414804 308218 414986 308454
rect 415222 308218 415404 308454
rect 414804 308134 415404 308218
rect 414804 307898 414986 308134
rect 415222 307898 415404 308134
rect 414804 274600 415404 307898
rect 432804 362454 433404 382916
rect 432804 362218 432986 362454
rect 433222 362218 433404 362454
rect 432804 362134 433404 362218
rect 432804 361898 432986 362134
rect 433222 361898 433404 362134
rect 432804 326454 433404 361898
rect 432804 326218 432986 326454
rect 433222 326218 433404 326454
rect 432804 326134 433404 326218
rect 432804 325898 432986 326134
rect 433222 325898 433404 326134
rect 432804 290454 433404 325898
rect 432804 290218 432986 290454
rect 433222 290218 433404 290454
rect 432804 290134 433404 290218
rect 432804 289898 432986 290134
rect 433222 289898 433404 290134
rect 432804 274600 433404 289898
rect 450804 380454 451404 382916
rect 450804 380218 450986 380454
rect 451222 380218 451404 380454
rect 450804 380134 451404 380218
rect 450804 379898 450986 380134
rect 451222 379898 451404 380134
rect 450804 344454 451404 379898
rect 450804 344218 450986 344454
rect 451222 344218 451404 344454
rect 450804 344134 451404 344218
rect 450804 343898 450986 344134
rect 451222 343898 451404 344134
rect 450804 308454 451404 343898
rect 450804 308218 450986 308454
rect 451222 308218 451404 308454
rect 450804 308134 451404 308218
rect 450804 307898 450986 308134
rect 451222 307898 451404 308134
rect 450804 274600 451404 307898
rect 468804 362454 469404 382916
rect 468804 362218 468986 362454
rect 469222 362218 469404 362454
rect 468804 362134 469404 362218
rect 468804 361898 468986 362134
rect 469222 361898 469404 362134
rect 468804 326454 469404 361898
rect 468804 326218 468986 326454
rect 469222 326218 469404 326454
rect 468804 326134 469404 326218
rect 468804 325898 468986 326134
rect 469222 325898 469404 326134
rect 468804 290454 469404 325898
rect 468804 290218 468986 290454
rect 469222 290218 469404 290454
rect 468804 290134 469404 290218
rect 468804 289898 468986 290134
rect 469222 289898 469404 290134
rect 468804 274600 469404 289898
rect 486804 380454 487404 382916
rect 486804 380218 486986 380454
rect 487222 380218 487404 380454
rect 486804 380134 487404 380218
rect 486804 379898 486986 380134
rect 487222 379898 487404 380134
rect 486804 344454 487404 379898
rect 486804 344218 486986 344454
rect 487222 344218 487404 344454
rect 486804 344134 487404 344218
rect 486804 343898 486986 344134
rect 487222 343898 487404 344134
rect 486804 308454 487404 343898
rect 486804 308218 486986 308454
rect 487222 308218 487404 308454
rect 486804 308134 487404 308218
rect 486804 307898 486986 308134
rect 487222 307898 487404 308134
rect 486804 274600 487404 307898
rect 504804 362454 505404 382916
rect 504804 362218 504986 362454
rect 505222 362218 505404 362454
rect 504804 362134 505404 362218
rect 504804 361898 504986 362134
rect 505222 361898 505404 362134
rect 504804 326454 505404 361898
rect 504804 326218 504986 326454
rect 505222 326218 505404 326454
rect 504804 326134 505404 326218
rect 504804 325898 504986 326134
rect 505222 325898 505404 326134
rect 504804 290454 505404 325898
rect 504804 290218 504986 290454
rect 505222 290218 505404 290454
rect 504804 290134 505404 290218
rect 504804 289898 504986 290134
rect 505222 289898 505404 290134
rect 504804 274600 505404 289898
rect 522804 380454 523404 382916
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 274600 523404 307898
rect 540804 362454 541404 382916
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 274600 541404 289898
rect 558804 380454 559404 382916
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 274600 559404 307898
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 306419 272236 306485 272237
rect 306419 272172 306420 272236
rect 306484 272172 306485 272236
rect 306419 272171 306485 272172
rect 306804 272218 306986 272454
rect 307222 272218 307404 272454
rect 306804 272134 307404 272218
rect 306804 271898 306986 272134
rect 307222 271898 307404 272134
rect 306804 236454 307404 271898
rect 554256 254454 554576 254476
rect 554256 254218 554298 254454
rect 554534 254218 554576 254454
rect 554256 254134 554576 254218
rect 554256 253898 554298 254134
rect 554534 253898 554576 254134
rect 554256 253876 554576 253898
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 306804 236218 306986 236454
rect 307222 236218 307404 236454
rect 306804 236134 307404 236218
rect 306804 235898 306986 236134
rect 307222 235898 307404 236134
rect 306804 200454 307404 235898
rect 538896 236454 539216 236476
rect 538896 236218 538938 236454
rect 539174 236218 539216 236454
rect 538896 236134 539216 236218
rect 538896 235898 538938 236134
rect 539174 235898 539216 236134
rect 538896 235876 539216 235898
rect 554256 218454 554576 218476
rect 554256 218218 554298 218454
rect 554534 218218 554576 218454
rect 554256 218134 554576 218218
rect 554256 217898 554298 218134
rect 554534 217898 554576 218134
rect 554256 217876 554576 217898
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 306804 200218 306986 200454
rect 307222 200218 307404 200454
rect 306804 200134 307404 200218
rect 306804 199898 306986 200134
rect 307222 199898 307404 200134
rect 306804 164454 307404 199898
rect 538896 200454 539216 200476
rect 538896 200218 538938 200454
rect 539174 200218 539216 200454
rect 538896 200134 539216 200218
rect 538896 199898 538938 200134
rect 539174 199898 539216 200134
rect 538896 199876 539216 199898
rect 554256 182454 554576 182476
rect 554256 182218 554298 182454
rect 554534 182218 554576 182454
rect 554256 182134 554576 182218
rect 554256 181898 554298 182134
rect 554534 181898 554576 182134
rect 554256 181876 554576 181898
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 306804 164218 306986 164454
rect 307222 164218 307404 164454
rect 306804 164134 307404 164218
rect 306804 163898 306986 164134
rect 307222 163898 307404 164134
rect 306804 128454 307404 163898
rect 538896 164454 539216 164476
rect 538896 164218 538938 164454
rect 539174 164218 539216 164454
rect 538896 164134 539216 164218
rect 538896 163898 538938 164134
rect 539174 163898 539216 164134
rect 538896 163876 539216 163898
rect 554256 146454 554576 146476
rect 554256 146218 554298 146454
rect 554534 146218 554576 146454
rect 554256 146134 554576 146218
rect 554256 145898 554298 146134
rect 554534 145898 554576 146134
rect 554256 145876 554576 145898
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 306804 128218 306986 128454
rect 307222 128218 307404 128454
rect 306804 128134 307404 128218
rect 306804 127898 306986 128134
rect 307222 127898 307404 128134
rect 306804 92454 307404 127898
rect 538896 128454 539216 128476
rect 538896 128218 538938 128454
rect 539174 128218 539216 128454
rect 538896 128134 539216 128218
rect 538896 127898 538938 128134
rect 539174 127898 539216 128134
rect 538896 127876 539216 127898
rect 554256 110454 554576 110476
rect 554256 110218 554298 110454
rect 554534 110218 554576 110454
rect 554256 110134 554576 110218
rect 554256 109898 554298 110134
rect 554534 109898 554576 110134
rect 554256 109876 554576 109898
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 300899 72044 300965 72045
rect 300899 71980 300900 72044
rect 300964 71980 300965 72044
rect 300899 71979 300965 71980
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1864 289404 -902
rect 306804 56454 307404 91898
rect 538896 92454 539216 92476
rect 538896 92218 538938 92454
rect 539174 92218 539216 92454
rect 538896 92134 539216 92218
rect 538896 91898 538938 92134
rect 539174 91898 539216 92134
rect 538896 91876 539216 91898
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1286 307404 19898
rect 306804 -1522 306986 -1286
rect 307222 -1522 307404 -1286
rect 306804 -1606 307404 -1522
rect 306804 -1842 306986 -1606
rect 307222 -1842 307404 -1606
rect 306804 -1864 307404 -1842
rect 324804 38454 325404 72600
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1864 325404 -902
rect 342804 56454 343404 72600
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1286 343404 19898
rect 342804 -1522 342986 -1286
rect 343222 -1522 343404 -1286
rect 342804 -1606 343404 -1522
rect 342804 -1842 342986 -1606
rect 343222 -1842 343404 -1606
rect 342804 -1864 343404 -1842
rect 360804 38454 361404 72600
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1864 361404 -902
rect 378804 56454 379404 72600
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1286 379404 19898
rect 378804 -1522 378986 -1286
rect 379222 -1522 379404 -1286
rect 378804 -1606 379404 -1522
rect 378804 -1842 378986 -1606
rect 379222 -1842 379404 -1606
rect 378804 -1864 379404 -1842
rect 396804 38454 397404 72600
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1864 397404 -902
rect 414804 56454 415404 72600
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1286 415404 19898
rect 414804 -1522 414986 -1286
rect 415222 -1522 415404 -1286
rect 414804 -1606 415404 -1522
rect 414804 -1842 414986 -1606
rect 415222 -1842 415404 -1606
rect 414804 -1864 415404 -1842
rect 432804 38454 433404 72600
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1864 433404 -902
rect 450804 56454 451404 72600
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1286 451404 19898
rect 450804 -1522 450986 -1286
rect 451222 -1522 451404 -1286
rect 450804 -1606 451404 -1522
rect 450804 -1842 450986 -1606
rect 451222 -1842 451404 -1606
rect 450804 -1864 451404 -1842
rect 468804 38454 469404 72600
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1864 469404 -902
rect 486804 56454 487404 72600
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1286 487404 19898
rect 486804 -1522 486986 -1286
rect 487222 -1522 487404 -1286
rect 486804 -1606 487404 -1522
rect 486804 -1842 486986 -1606
rect 487222 -1842 487404 -1606
rect 486804 -1864 487404 -1842
rect 504804 38454 505404 72600
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1864 505404 -902
rect 522804 56454 523404 72600
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1286 523404 19898
rect 522804 -1522 522986 -1286
rect 523222 -1522 523404 -1286
rect 522804 -1606 523404 -1522
rect 522804 -1842 522986 -1606
rect 523222 -1842 523404 -1606
rect 522804 -1864 523404 -1842
rect 540804 38454 541404 72600
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1864 541404 -902
rect 558804 56454 559404 72600
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1286 559404 19898
rect 558804 -1522 558986 -1286
rect 559222 -1522 559404 -1286
rect 558804 -1606 559404 -1522
rect 558804 -1842 558986 -1606
rect 559222 -1842 559404 -1606
rect 558804 -1864 559404 -1842
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1864 577404 -902
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586260 668454 586860 705222
rect 586260 668218 586442 668454
rect 586678 668218 586860 668454
rect 586260 668134 586860 668218
rect 586260 667898 586442 668134
rect 586678 667898 586860 668134
rect 586260 632454 586860 667898
rect 586260 632218 586442 632454
rect 586678 632218 586860 632454
rect 586260 632134 586860 632218
rect 586260 631898 586442 632134
rect 586678 631898 586860 632134
rect 586260 596454 586860 631898
rect 586260 596218 586442 596454
rect 586678 596218 586860 596454
rect 586260 596134 586860 596218
rect 586260 595898 586442 596134
rect 586678 595898 586860 596134
rect 586260 560454 586860 595898
rect 586260 560218 586442 560454
rect 586678 560218 586860 560454
rect 586260 560134 586860 560218
rect 586260 559898 586442 560134
rect 586678 559898 586860 560134
rect 586260 524454 586860 559898
rect 586260 524218 586442 524454
rect 586678 524218 586860 524454
rect 586260 524134 586860 524218
rect 586260 523898 586442 524134
rect 586678 523898 586860 524134
rect 586260 488454 586860 523898
rect 586260 488218 586442 488454
rect 586678 488218 586860 488454
rect 586260 488134 586860 488218
rect 586260 487898 586442 488134
rect 586678 487898 586860 488134
rect 586260 452454 586860 487898
rect 586260 452218 586442 452454
rect 586678 452218 586860 452454
rect 586260 452134 586860 452218
rect 586260 451898 586442 452134
rect 586678 451898 586860 452134
rect 586260 416454 586860 451898
rect 586260 416218 586442 416454
rect 586678 416218 586860 416454
rect 586260 416134 586860 416218
rect 586260 415898 586442 416134
rect 586678 415898 586860 416134
rect 586260 380454 586860 415898
rect 586260 380218 586442 380454
rect 586678 380218 586860 380454
rect 586260 380134 586860 380218
rect 586260 379898 586442 380134
rect 586678 379898 586860 380134
rect 586260 344454 586860 379898
rect 586260 344218 586442 344454
rect 586678 344218 586860 344454
rect 586260 344134 586860 344218
rect 586260 343898 586442 344134
rect 586678 343898 586860 344134
rect 586260 308454 586860 343898
rect 586260 308218 586442 308454
rect 586678 308218 586860 308454
rect 586260 308134 586860 308218
rect 586260 307898 586442 308134
rect 586678 307898 586860 308134
rect 586260 272454 586860 307898
rect 586260 272218 586442 272454
rect 586678 272218 586860 272454
rect 586260 272134 586860 272218
rect 586260 271898 586442 272134
rect 586678 271898 586860 272134
rect 586260 236454 586860 271898
rect 586260 236218 586442 236454
rect 586678 236218 586860 236454
rect 586260 236134 586860 236218
rect 586260 235898 586442 236134
rect 586678 235898 586860 236134
rect 586260 200454 586860 235898
rect 586260 200218 586442 200454
rect 586678 200218 586860 200454
rect 586260 200134 586860 200218
rect 586260 199898 586442 200134
rect 586678 199898 586860 200134
rect 586260 164454 586860 199898
rect 586260 164218 586442 164454
rect 586678 164218 586860 164454
rect 586260 164134 586860 164218
rect 586260 163898 586442 164134
rect 586678 163898 586860 164134
rect 586260 128454 586860 163898
rect 586260 128218 586442 128454
rect 586678 128218 586860 128454
rect 586260 128134 586860 128218
rect 586260 127898 586442 128134
rect 586678 127898 586860 128134
rect 586260 92454 586860 127898
rect 586260 92218 586442 92454
rect 586678 92218 586860 92454
rect 586260 92134 586860 92218
rect 586260 91898 586442 92134
rect 586678 91898 586860 92134
rect 586260 56454 586860 91898
rect 586260 56218 586442 56454
rect 586678 56218 586860 56454
rect 586260 56134 586860 56218
rect 586260 55898 586442 56134
rect 586678 55898 586860 56134
rect 586260 20454 586860 55898
rect 586260 20218 586442 20454
rect 586678 20218 586860 20454
rect 586260 20134 586860 20218
rect 586260 19898 586442 20134
rect 586678 19898 586860 20134
rect 586260 -1286 586860 19898
rect 586260 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect 586260 -1606 586860 -1522
rect 586260 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect 586260 -1864 586860 -1842
rect -3876 -2462 -3694 -2226
rect -3458 -2462 -3276 -2226
rect -3876 -2546 -3276 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 -3276 -2546
rect -3876 -2804 -3276 -2782
rect 587200 -2226 587800 706162
rect 587200 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect 587200 -2546 587800 -2462
rect 587200 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect 587200 -2804 587800 -2782
rect -4816 -3402 -4634 -3166
rect -4398 -3402 -4216 -3166
rect -4816 -3486 -4216 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 -4216 -3486
rect -4816 -3744 -4216 -3722
rect 588140 -3166 588740 707102
rect 588140 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect 588140 -3486 588740 -3402
rect 588140 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect 588140 -3744 588740 -3722
rect -5756 -4342 -5574 -4106
rect -5338 -4342 -5156 -4106
rect -5756 -4426 -5156 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 -5156 -4426
rect -5756 -4684 -5156 -4662
rect 589080 -4106 589680 708042
rect 589080 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect 589080 -4426 589680 -4342
rect 589080 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect 589080 -4684 589680 -4662
rect -6696 -5282 -6514 -5046
rect -6278 -5282 -6096 -5046
rect -6696 -5366 -6096 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 -6096 -5366
rect -6696 -5624 -6096 -5602
rect 590020 -5046 590620 708982
rect 590020 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect 590020 -5366 590620 -5282
rect 590020 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect 590020 -5624 590620 -5602
rect -7636 -6222 -7454 -5986
rect -7218 -6222 -7036 -5986
rect -7636 -6306 -7036 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 -7036 -6306
rect -7636 -6564 -7036 -6542
rect 590960 -5986 591560 709922
rect 590960 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect 590960 -6306 591560 -6222
rect 590960 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect 590960 -6564 591560 -6542
rect -8576 -7162 -8394 -6926
rect -8158 -7162 -7976 -6926
rect -8576 -7246 -7976 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 -7976 -7246
rect -8576 -7504 -7976 -7482
rect 591900 -6926 592500 710862
rect 591900 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect 591900 -7246 592500 -7162
rect 591900 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect 591900 -7504 592500 -7482
<< via4 >>
rect -8394 711182 -8158 711418
rect -8394 710862 -8158 711098
rect 592082 711182 592318 711418
rect 592082 710862 592318 711098
rect -7454 710242 -7218 710478
rect -7454 709922 -7218 710158
rect 591142 710242 591378 710478
rect 591142 709922 591378 710158
rect -6514 709302 -6278 709538
rect -6514 708982 -6278 709218
rect 590202 709302 590438 709538
rect 590202 708982 590438 709218
rect -5574 708362 -5338 708598
rect -5574 708042 -5338 708278
rect 589262 708362 589498 708598
rect 589262 708042 589498 708278
rect -4634 707422 -4398 707658
rect -4634 707102 -4398 707338
rect 588322 707422 588558 707658
rect 588322 707102 588558 707338
rect -3694 706482 -3458 706718
rect -3694 706162 -3458 706398
rect 587382 706482 587618 706718
rect 587382 706162 587618 706398
rect -2754 705542 -2518 705778
rect -2754 705222 -2518 705458
rect -2754 668218 -2518 668454
rect -2754 667898 -2518 668134
rect -2754 632218 -2518 632454
rect -2754 631898 -2518 632134
rect -2754 596218 -2518 596454
rect -2754 595898 -2518 596134
rect -2754 560218 -2518 560454
rect -2754 559898 -2518 560134
rect -2754 524218 -2518 524454
rect -2754 523898 -2518 524134
rect -2754 488218 -2518 488454
rect -2754 487898 -2518 488134
rect -2754 452218 -2518 452454
rect -2754 451898 -2518 452134
rect -2754 416218 -2518 416454
rect -2754 415898 -2518 416134
rect -2754 380218 -2518 380454
rect -2754 379898 -2518 380134
rect -2754 344218 -2518 344454
rect -2754 343898 -2518 344134
rect -2754 308218 -2518 308454
rect -2754 307898 -2518 308134
rect -2754 272218 -2518 272454
rect -2754 271898 -2518 272134
rect -2754 236218 -2518 236454
rect -2754 235898 -2518 236134
rect -2754 200218 -2518 200454
rect -2754 199898 -2518 200134
rect -2754 164218 -2518 164454
rect -2754 163898 -2518 164134
rect -2754 128218 -2518 128454
rect -2754 127898 -2518 128134
rect -2754 92218 -2518 92454
rect -2754 91898 -2518 92134
rect -2754 56218 -2518 56454
rect -2754 55898 -2518 56134
rect -2754 20218 -2518 20454
rect -2754 19898 -2518 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2754 -1522 -2518 -1286
rect -2754 -1842 -2518 -1606
rect 18986 705542 19222 705778
rect 18986 705222 19222 705458
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 54986 705542 55222 705778
rect 54986 705222 55222 705458
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 72986 614218 73222 614454
rect 72986 613898 73222 614134
rect 90986 705542 91222 705778
rect 90986 705222 91222 705458
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 90986 632218 91222 632454
rect 90986 631898 91222 632134
rect 90986 596218 91222 596454
rect 90986 595898 91222 596134
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 108986 614218 109222 614454
rect 108986 613898 109222 614134
rect 126986 705542 127222 705778
rect 126986 705222 127222 705458
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 126986 632218 127222 632454
rect 126986 631898 127222 632134
rect 126986 596218 127222 596454
rect 126986 595898 127222 596134
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 162986 705542 163222 705778
rect 162986 705222 163222 705458
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 198986 705542 199222 705778
rect 198986 705222 199222 705458
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 198986 632218 199222 632454
rect 198986 631898 199222 632134
rect 198986 596218 199222 596454
rect 198986 595898 199222 596134
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 216986 614218 217222 614454
rect 216986 613898 217222 614134
rect 234986 705542 235222 705778
rect 234986 705222 235222 705458
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 234986 632218 235222 632454
rect 234986 631898 235222 632134
rect 234986 596218 235222 596454
rect 234986 595898 235222 596134
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 252986 614218 253222 614454
rect 252986 613898 253222 614134
rect 270986 705542 271222 705778
rect 270986 705222 271222 705458
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 270986 596218 271222 596454
rect 270986 595898 271222 596134
rect 262170 578218 262406 578454
rect 262170 577898 262406 578134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 246810 560218 247046 560454
rect 246810 559898 247046 560134
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 262170 542218 262406 542454
rect 262170 541898 262406 542134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 246810 524218 247046 524454
rect 246810 523898 247046 524134
rect 270986 524218 271222 524454
rect 270986 523898 271222 524134
rect 262170 506218 262406 506454
rect 262170 505898 262406 506134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 246810 488218 247046 488454
rect 246810 487898 247046 488134
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 306986 705542 307222 705778
rect 306986 705222 307222 705458
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 306986 596218 307222 596454
rect 306986 595898 307222 596134
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 288986 542218 289222 542454
rect 288986 541898 289222 542134
rect 270986 488218 271222 488454
rect 270986 487898 271222 488134
rect 262170 470218 262406 470454
rect 262170 469898 262406 470134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 246810 452218 247046 452454
rect 246810 451898 247046 452134
rect 270986 452218 271222 452454
rect 270986 451898 271222 452134
rect 262170 434218 262406 434454
rect 262170 433898 262406 434134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 246810 416218 247046 416454
rect 246810 415898 247046 416134
rect 270986 416218 271222 416454
rect 270986 415898 271222 416134
rect 262170 398218 262406 398454
rect 262170 397898 262406 398134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 72986 362218 73222 362454
rect 72986 361898 73222 362134
rect 72986 326218 73222 326454
rect 72986 325898 73222 326134
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 90986 380218 91222 380454
rect 90986 379898 91222 380134
rect 90986 344218 91222 344454
rect 90986 343898 91222 344134
rect 90986 308218 91222 308454
rect 90986 307898 91222 308134
rect 108986 362218 109222 362454
rect 108986 361898 109222 362134
rect 108986 326218 109222 326454
rect 108986 325898 109222 326134
rect 108986 290218 109222 290454
rect 108986 289898 109222 290134
rect 126986 380218 127222 380454
rect 126986 379898 127222 380134
rect 126986 344218 127222 344454
rect 126986 343898 127222 344134
rect 126986 308218 127222 308454
rect 126986 307898 127222 308134
rect 144986 362218 145222 362454
rect 144986 361898 145222 362134
rect 144986 326218 145222 326454
rect 144986 325898 145222 326134
rect 144986 290218 145222 290454
rect 144986 289898 145222 290134
rect 162986 380218 163222 380454
rect 162986 379898 163222 380134
rect 162986 344218 163222 344454
rect 162986 343898 163222 344134
rect 162986 308218 163222 308454
rect 162986 307898 163222 308134
rect 180986 362218 181222 362454
rect 180986 361898 181222 362134
rect 180986 326218 181222 326454
rect 180986 325898 181222 326134
rect 180986 290218 181222 290454
rect 180986 289898 181222 290134
rect 198986 380218 199222 380454
rect 198986 379898 199222 380134
rect 198986 344218 199222 344454
rect 198986 343898 199222 344134
rect 198986 308218 199222 308454
rect 198986 307898 199222 308134
rect 216986 362218 217222 362454
rect 216986 361898 217222 362134
rect 216986 326218 217222 326454
rect 216986 325898 217222 326134
rect 216986 290218 217222 290454
rect 216986 289898 217222 290134
rect 234986 380218 235222 380454
rect 234986 379898 235222 380134
rect 234986 344218 235222 344454
rect 234986 343898 235222 344134
rect 234986 308218 235222 308454
rect 234986 307898 235222 308134
rect 252986 362218 253222 362454
rect 252986 361898 253222 362134
rect 270986 380218 271222 380454
rect 270986 379898 271222 380134
rect 252986 326218 253222 326454
rect 252986 325898 253222 326134
rect 252986 290218 253222 290454
rect 252986 289898 253222 290134
rect 270986 308218 271222 308454
rect 270986 307898 271222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 288986 506218 289222 506454
rect 288986 505898 289222 506134
rect 288986 470218 289222 470454
rect 288986 469898 289222 470134
rect 288986 434218 289222 434454
rect 288986 433898 289222 434134
rect 288986 398218 289222 398454
rect 288986 397898 289222 398134
rect 288986 362218 289222 362454
rect 288986 361898 289222 362134
rect 270986 272218 271222 272454
rect 270986 271898 271222 272134
rect 262170 254218 262406 254454
rect 262170 253898 262406 254134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 246810 236218 247046 236454
rect 246810 235898 247046 236134
rect 270986 236218 271222 236454
rect 270986 235898 271222 236134
rect 262170 218218 262406 218454
rect 262170 217898 262406 218134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 246810 200218 247046 200454
rect 246810 199898 247046 200134
rect 270986 200218 271222 200454
rect 270986 199898 271222 200134
rect 262170 182218 262406 182454
rect 262170 181898 262406 182134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 246810 164218 247046 164454
rect 246810 163898 247046 164134
rect 270986 164218 271222 164454
rect 270986 163898 271222 164134
rect 262170 146218 262406 146454
rect 262170 145898 262406 146134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 246810 128218 247046 128454
rect 246810 127898 247046 128134
rect 270986 128218 271222 128454
rect 270986 127898 271222 128134
rect 262170 110218 262406 110454
rect 262170 109898 262406 110134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 246810 92218 247046 92454
rect 246810 91898 247046 92134
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1522 19222 -1286
rect 18986 -1842 19222 -1606
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1522 55222 -1286
rect 54986 -1842 55222 -1606
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1522 91222 -1286
rect 90986 -1842 91222 -1606
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1522 127222 -1286
rect 126986 -1842 127222 -1606
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1522 163222 -1286
rect 162986 -1842 163222 -1606
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1522 199222 -1286
rect 198986 -1842 199222 -1606
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1522 235222 -1286
rect 234986 -1842 235222 -1606
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 288986 290218 289222 290454
rect 288986 289898 289222 290134
rect 292154 344218 292390 344454
rect 292154 343898 292390 344134
rect 288986 254218 289222 254454
rect 288986 253898 289222 254134
rect 288986 218218 289222 218454
rect 288986 217898 289222 218134
rect 288986 182218 289222 182454
rect 288986 181898 289222 182134
rect 288986 146218 289222 146454
rect 288986 145898 289222 146134
rect 288986 110218 289222 110454
rect 288986 109898 289222 110134
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1522 271222 -1286
rect 270986 -1842 271222 -1606
rect 306986 560218 307222 560454
rect 306986 559898 307222 560134
rect 306986 524218 307222 524454
rect 306986 523898 307222 524134
rect 306986 488218 307222 488454
rect 306986 487898 307222 488134
rect 306986 452218 307222 452454
rect 306986 451898 307222 452134
rect 306986 416218 307222 416454
rect 306986 415898 307222 416134
rect 306986 380218 307222 380454
rect 306986 379898 307222 380134
rect 307514 326218 307750 326454
rect 307514 325898 307750 326134
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 324986 650218 325222 650454
rect 324986 649898 325222 650134
rect 324986 614218 325222 614454
rect 324986 613898 325222 614134
rect 342986 705542 343222 705778
rect 342986 705222 343222 705458
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 342986 632218 343222 632454
rect 342986 631898 343222 632134
rect 342986 596218 343222 596454
rect 342986 595898 343222 596134
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 360986 650218 361222 650454
rect 360986 649898 361222 650134
rect 360986 614218 361222 614454
rect 360986 613898 361222 614134
rect 378986 705542 379222 705778
rect 378986 705222 379222 705458
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 378986 632218 379222 632454
rect 378986 631898 379222 632134
rect 378986 596218 379222 596454
rect 378986 595898 379222 596134
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 414986 705542 415222 705778
rect 414986 705222 415222 705458
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 414986 596218 415222 596454
rect 414986 595898 415222 596134
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 450986 705542 451222 705778
rect 450986 705222 451222 705458
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 450986 632218 451222 632454
rect 450986 631898 451222 632134
rect 450986 596218 451222 596454
rect 450986 595898 451222 596134
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 468986 614218 469222 614454
rect 468986 613898 469222 614134
rect 486986 705542 487222 705778
rect 486986 705222 487222 705458
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 486986 632218 487222 632454
rect 486986 631898 487222 632134
rect 486986 596218 487222 596454
rect 486986 595898 487222 596134
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 504986 614218 505222 614454
rect 504986 613898 505222 614134
rect 522986 705542 523222 705778
rect 522986 705222 523222 705458
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 558986 705542 559222 705778
rect 558986 705222 559222 705458
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 586442 705542 586678 705778
rect 586442 705222 586678 705458
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 554298 578218 554534 578454
rect 554298 577898 554534 578134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 538938 560218 539174 560454
rect 538938 559898 539174 560134
rect 554298 542218 554534 542454
rect 554298 541898 554534 542134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 538938 524218 539174 524454
rect 538938 523898 539174 524134
rect 554298 506218 554534 506454
rect 554298 505898 554534 506134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 538938 488218 539174 488454
rect 538938 487898 539174 488134
rect 554298 470218 554534 470454
rect 554298 469898 554534 470134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 538938 452218 539174 452454
rect 538938 451898 539174 452134
rect 554298 434218 554534 434454
rect 554298 433898 554534 434134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 538938 416218 539174 416454
rect 538938 415898 539174 416134
rect 554298 398218 554534 398454
rect 554298 397898 554534 398134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 324986 362218 325222 362454
rect 324986 361898 325222 362134
rect 324986 326218 325222 326454
rect 324986 325898 325222 326134
rect 306986 308218 307222 308454
rect 306986 307898 307222 308134
rect 324986 290218 325222 290454
rect 324986 289898 325222 290134
rect 342986 380218 343222 380454
rect 342986 379898 343222 380134
rect 342986 344218 343222 344454
rect 342986 343898 343222 344134
rect 342986 308218 343222 308454
rect 342986 307898 343222 308134
rect 360986 362218 361222 362454
rect 360986 361898 361222 362134
rect 360986 326218 361222 326454
rect 360986 325898 361222 326134
rect 360986 290218 361222 290454
rect 360986 289898 361222 290134
rect 378986 380218 379222 380454
rect 378986 379898 379222 380134
rect 378986 344218 379222 344454
rect 378986 343898 379222 344134
rect 378986 308218 379222 308454
rect 378986 307898 379222 308134
rect 396986 362218 397222 362454
rect 396986 361898 397222 362134
rect 396986 326218 397222 326454
rect 396986 325898 397222 326134
rect 396986 290218 397222 290454
rect 396986 289898 397222 290134
rect 414986 380218 415222 380454
rect 414986 379898 415222 380134
rect 414986 344218 415222 344454
rect 414986 343898 415222 344134
rect 414986 308218 415222 308454
rect 414986 307898 415222 308134
rect 432986 362218 433222 362454
rect 432986 361898 433222 362134
rect 432986 326218 433222 326454
rect 432986 325898 433222 326134
rect 432986 290218 433222 290454
rect 432986 289898 433222 290134
rect 450986 380218 451222 380454
rect 450986 379898 451222 380134
rect 450986 344218 451222 344454
rect 450986 343898 451222 344134
rect 450986 308218 451222 308454
rect 450986 307898 451222 308134
rect 468986 362218 469222 362454
rect 468986 361898 469222 362134
rect 468986 326218 469222 326454
rect 468986 325898 469222 326134
rect 468986 290218 469222 290454
rect 468986 289898 469222 290134
rect 486986 380218 487222 380454
rect 486986 379898 487222 380134
rect 486986 344218 487222 344454
rect 486986 343898 487222 344134
rect 486986 308218 487222 308454
rect 486986 307898 487222 308134
rect 504986 362218 505222 362454
rect 504986 361898 505222 362134
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 306986 272218 307222 272454
rect 306986 271898 307222 272134
rect 554298 254218 554534 254454
rect 554298 253898 554534 254134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 306986 236218 307222 236454
rect 306986 235898 307222 236134
rect 538938 236218 539174 236454
rect 538938 235898 539174 236134
rect 554298 218218 554534 218454
rect 554298 217898 554534 218134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 306986 200218 307222 200454
rect 306986 199898 307222 200134
rect 538938 200218 539174 200454
rect 538938 199898 539174 200134
rect 554298 182218 554534 182454
rect 554298 181898 554534 182134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 306986 164218 307222 164454
rect 306986 163898 307222 164134
rect 538938 164218 539174 164454
rect 538938 163898 539174 164134
rect 554298 146218 554534 146454
rect 554298 145898 554534 146134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 306986 128218 307222 128454
rect 306986 127898 307222 128134
rect 538938 128218 539174 128454
rect 538938 127898 539174 128134
rect 554298 110218 554534 110454
rect 554298 109898 554534 110134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 538938 92218 539174 92454
rect 538938 91898 539174 92134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1522 307222 -1286
rect 306986 -1842 307222 -1606
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1522 343222 -1286
rect 342986 -1842 343222 -1606
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1522 379222 -1286
rect 378986 -1842 379222 -1606
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1522 415222 -1286
rect 414986 -1842 415222 -1606
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1522 451222 -1286
rect 450986 -1842 451222 -1606
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1522 487222 -1286
rect 486986 -1842 487222 -1606
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1522 523222 -1286
rect 522986 -1842 523222 -1606
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1522 559222 -1286
rect 558986 -1842 559222 -1606
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586442 668218 586678 668454
rect 586442 667898 586678 668134
rect 586442 632218 586678 632454
rect 586442 631898 586678 632134
rect 586442 596218 586678 596454
rect 586442 595898 586678 596134
rect 586442 560218 586678 560454
rect 586442 559898 586678 560134
rect 586442 524218 586678 524454
rect 586442 523898 586678 524134
rect 586442 488218 586678 488454
rect 586442 487898 586678 488134
rect 586442 452218 586678 452454
rect 586442 451898 586678 452134
rect 586442 416218 586678 416454
rect 586442 415898 586678 416134
rect 586442 380218 586678 380454
rect 586442 379898 586678 380134
rect 586442 344218 586678 344454
rect 586442 343898 586678 344134
rect 586442 308218 586678 308454
rect 586442 307898 586678 308134
rect 586442 272218 586678 272454
rect 586442 271898 586678 272134
rect 586442 236218 586678 236454
rect 586442 235898 586678 236134
rect 586442 200218 586678 200454
rect 586442 199898 586678 200134
rect 586442 164218 586678 164454
rect 586442 163898 586678 164134
rect 586442 128218 586678 128454
rect 586442 127898 586678 128134
rect 586442 92218 586678 92454
rect 586442 91898 586678 92134
rect 586442 56218 586678 56454
rect 586442 55898 586678 56134
rect 586442 20218 586678 20454
rect 586442 19898 586678 20134
rect 586442 -1522 586678 -1286
rect 586442 -1842 586678 -1606
rect -3694 -2462 -3458 -2226
rect -3694 -2782 -3458 -2546
rect 587382 -2462 587618 -2226
rect 587382 -2782 587618 -2546
rect -4634 -3402 -4398 -3166
rect -4634 -3722 -4398 -3486
rect 588322 -3402 588558 -3166
rect 588322 -3722 588558 -3486
rect -5574 -4342 -5338 -4106
rect -5574 -4662 -5338 -4426
rect 589262 -4342 589498 -4106
rect 589262 -4662 589498 -4426
rect -6514 -5282 -6278 -5046
rect -6514 -5602 -6278 -5366
rect 590202 -5282 590438 -5046
rect 590202 -5602 590438 -5366
rect -7454 -6222 -7218 -5986
rect -7454 -6542 -7218 -6306
rect 591142 -6222 591378 -5986
rect 591142 -6542 591378 -6306
rect -8394 -7162 -8158 -6926
rect -8394 -7482 -8158 -7246
rect 592082 -7162 592318 -6926
rect 592082 -7482 592318 -7246
<< metal5 >>
rect -8576 711440 -7976 711442
rect 591900 711440 592500 711442
rect -8576 711418 592500 711440
rect -8576 711182 -8394 711418
rect -8158 711182 592082 711418
rect 592318 711182 592500 711418
rect -8576 711098 592500 711182
rect -8576 710862 -8394 711098
rect -8158 710862 592082 711098
rect 592318 710862 592500 711098
rect -8576 710840 592500 710862
rect -8576 710838 -7976 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 590960 710500 591560 710502
rect -7636 710478 591560 710500
rect -7636 710242 -7454 710478
rect -7218 710242 591142 710478
rect 591378 710242 591560 710478
rect -7636 710158 591560 710242
rect -7636 709922 -7454 710158
rect -7218 709922 591142 710158
rect 591378 709922 591560 710158
rect -7636 709900 591560 709922
rect -7636 709898 -7036 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 590020 709560 590620 709562
rect -6696 709538 590620 709560
rect -6696 709302 -6514 709538
rect -6278 709302 590202 709538
rect 590438 709302 590620 709538
rect -6696 709218 590620 709302
rect -6696 708982 -6514 709218
rect -6278 708982 590202 709218
rect 590438 708982 590620 709218
rect -6696 708960 590620 708982
rect -6696 708958 -6096 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 589080 708620 589680 708622
rect -5756 708598 589680 708620
rect -5756 708362 -5574 708598
rect -5338 708362 589262 708598
rect 589498 708362 589680 708598
rect -5756 708278 589680 708362
rect -5756 708042 -5574 708278
rect -5338 708042 589262 708278
rect 589498 708042 589680 708278
rect -5756 708020 589680 708042
rect -5756 708018 -5156 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 588140 707680 588740 707682
rect -4816 707658 588740 707680
rect -4816 707422 -4634 707658
rect -4398 707422 588322 707658
rect 588558 707422 588740 707658
rect -4816 707338 588740 707422
rect -4816 707102 -4634 707338
rect -4398 707102 588322 707338
rect 588558 707102 588740 707338
rect -4816 707080 588740 707102
rect -4816 707078 -4216 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 587200 706740 587800 706742
rect -3876 706718 587800 706740
rect -3876 706482 -3694 706718
rect -3458 706482 587382 706718
rect 587618 706482 587800 706718
rect -3876 706398 587800 706482
rect -3876 706162 -3694 706398
rect -3458 706162 587382 706398
rect 587618 706162 587800 706398
rect -3876 706140 587800 706162
rect -3876 706138 -3276 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 18804 705800 19404 705802
rect 54804 705800 55404 705802
rect 90804 705800 91404 705802
rect 126804 705800 127404 705802
rect 162804 705800 163404 705802
rect 198804 705800 199404 705802
rect 234804 705800 235404 705802
rect 270804 705800 271404 705802
rect 306804 705800 307404 705802
rect 342804 705800 343404 705802
rect 378804 705800 379404 705802
rect 414804 705800 415404 705802
rect 450804 705800 451404 705802
rect 486804 705800 487404 705802
rect 522804 705800 523404 705802
rect 558804 705800 559404 705802
rect 586260 705800 586860 705802
rect -2936 705778 586860 705800
rect -2936 705542 -2754 705778
rect -2518 705542 18986 705778
rect 19222 705542 54986 705778
rect 55222 705542 90986 705778
rect 91222 705542 126986 705778
rect 127222 705542 162986 705778
rect 163222 705542 198986 705778
rect 199222 705542 234986 705778
rect 235222 705542 270986 705778
rect 271222 705542 306986 705778
rect 307222 705542 342986 705778
rect 343222 705542 378986 705778
rect 379222 705542 414986 705778
rect 415222 705542 450986 705778
rect 451222 705542 486986 705778
rect 487222 705542 522986 705778
rect 523222 705542 558986 705778
rect 559222 705542 586442 705778
rect 586678 705542 586860 705778
rect -2936 705458 586860 705542
rect -2936 705222 -2754 705458
rect -2518 705222 18986 705458
rect 19222 705222 54986 705458
rect 55222 705222 90986 705458
rect 91222 705222 126986 705458
rect 127222 705222 162986 705458
rect 163222 705222 198986 705458
rect 199222 705222 234986 705458
rect 235222 705222 270986 705458
rect 271222 705222 306986 705458
rect 307222 705222 342986 705458
rect 343222 705222 378986 705458
rect 379222 705222 414986 705458
rect 415222 705222 450986 705458
rect 451222 705222 486986 705458
rect 487222 705222 522986 705458
rect 523222 705222 558986 705458
rect 559222 705222 586442 705458
rect 586678 705222 586860 705458
rect -2936 705200 586860 705222
rect -2936 705198 -2336 705200
rect 18804 705198 19404 705200
rect 54804 705198 55404 705200
rect 90804 705198 91404 705200
rect 126804 705198 127404 705200
rect 162804 705198 163404 705200
rect 198804 705198 199404 705200
rect 234804 705198 235404 705200
rect 270804 705198 271404 705200
rect 306804 705198 307404 705200
rect 342804 705198 343404 705200
rect 378804 705198 379404 705200
rect 414804 705198 415404 705200
rect 450804 705198 451404 705200
rect 486804 705198 487404 705200
rect 522804 705198 523404 705200
rect 558804 705198 559404 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2936 686454 586860 686476
rect -2936 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586860 686454
rect -2936 686134 586860 686218
rect -2936 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586860 686134
rect -2936 685876 586860 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -2936 668476 -2336 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586260 668476 586860 668478
rect -2936 668454 586860 668476
rect -2936 668218 -2754 668454
rect -2518 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586442 668454
rect 586678 668218 586860 668454
rect -2936 668134 586860 668218
rect -2936 667898 -2754 668134
rect -2518 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586442 668134
rect 586678 667898 586860 668134
rect -2936 667876 586860 667898
rect -2936 667874 -2336 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586260 667874 586860 667876
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 108804 650476 109404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 216804 650476 217404 650478
rect 252804 650476 253404 650478
rect 288804 650476 289404 650478
rect 324804 650476 325404 650478
rect 360804 650476 361404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 468804 650476 469404 650478
rect 504804 650476 505404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2936 650454 586860 650476
rect -2936 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 324986 650454
rect 325222 650218 360986 650454
rect 361222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586860 650454
rect -2936 650134 586860 650218
rect -2936 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 324986 650134
rect 325222 649898 360986 650134
rect 361222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586860 650134
rect -2936 649876 586860 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 108804 649874 109404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 216804 649874 217404 649876
rect 252804 649874 253404 649876
rect 288804 649874 289404 649876
rect 324804 649874 325404 649876
rect 360804 649874 361404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 468804 649874 469404 649876
rect 504804 649874 505404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -2936 632476 -2336 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 90804 632476 91404 632478
rect 126804 632476 127404 632478
rect 162804 632476 163404 632478
rect 198804 632476 199404 632478
rect 234804 632476 235404 632478
rect 270804 632476 271404 632478
rect 306804 632476 307404 632478
rect 342804 632476 343404 632478
rect 378804 632476 379404 632478
rect 414804 632476 415404 632478
rect 450804 632476 451404 632478
rect 486804 632476 487404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586260 632476 586860 632478
rect -2936 632454 586860 632476
rect -2936 632218 -2754 632454
rect -2518 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 90986 632454
rect 91222 632218 126986 632454
rect 127222 632218 162986 632454
rect 163222 632218 198986 632454
rect 199222 632218 234986 632454
rect 235222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 342986 632454
rect 343222 632218 378986 632454
rect 379222 632218 414986 632454
rect 415222 632218 450986 632454
rect 451222 632218 486986 632454
rect 487222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586442 632454
rect 586678 632218 586860 632454
rect -2936 632134 586860 632218
rect -2936 631898 -2754 632134
rect -2518 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 90986 632134
rect 91222 631898 126986 632134
rect 127222 631898 162986 632134
rect 163222 631898 198986 632134
rect 199222 631898 234986 632134
rect 235222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 342986 632134
rect 343222 631898 378986 632134
rect 379222 631898 414986 632134
rect 415222 631898 450986 632134
rect 451222 631898 486986 632134
rect 487222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586442 632134
rect 586678 631898 586860 632134
rect -2936 631876 586860 631898
rect -2936 631874 -2336 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 90804 631874 91404 631876
rect 126804 631874 127404 631876
rect 162804 631874 163404 631876
rect 198804 631874 199404 631876
rect 234804 631874 235404 631876
rect 270804 631874 271404 631876
rect 306804 631874 307404 631876
rect 342804 631874 343404 631876
rect 378804 631874 379404 631876
rect 414804 631874 415404 631876
rect 450804 631874 451404 631876
rect 486804 631874 487404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586260 631874 586860 631876
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 72804 614476 73404 614478
rect 108804 614476 109404 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 216804 614476 217404 614478
rect 252804 614476 253404 614478
rect 288804 614476 289404 614478
rect 324804 614476 325404 614478
rect 360804 614476 361404 614478
rect 396804 614476 397404 614478
rect 432804 614476 433404 614478
rect 468804 614476 469404 614478
rect 504804 614476 505404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2936 614454 586860 614476
rect -2936 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 72986 614454
rect 73222 614218 108986 614454
rect 109222 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 216986 614454
rect 217222 614218 252986 614454
rect 253222 614218 288986 614454
rect 289222 614218 324986 614454
rect 325222 614218 360986 614454
rect 361222 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 468986 614454
rect 469222 614218 504986 614454
rect 505222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586860 614454
rect -2936 614134 586860 614218
rect -2936 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 72986 614134
rect 73222 613898 108986 614134
rect 109222 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 216986 614134
rect 217222 613898 252986 614134
rect 253222 613898 288986 614134
rect 289222 613898 324986 614134
rect 325222 613898 360986 614134
rect 361222 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 468986 614134
rect 469222 613898 504986 614134
rect 505222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586860 614134
rect -2936 613876 586860 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 72804 613874 73404 613876
rect 108804 613874 109404 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 216804 613874 217404 613876
rect 252804 613874 253404 613876
rect 288804 613874 289404 613876
rect 324804 613874 325404 613876
rect 360804 613874 361404 613876
rect 396804 613874 397404 613876
rect 432804 613874 433404 613876
rect 468804 613874 469404 613876
rect 504804 613874 505404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -2936 596476 -2336 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 90804 596476 91404 596478
rect 126804 596476 127404 596478
rect 162804 596476 163404 596478
rect 198804 596476 199404 596478
rect 234804 596476 235404 596478
rect 270804 596476 271404 596478
rect 306804 596476 307404 596478
rect 342804 596476 343404 596478
rect 378804 596476 379404 596478
rect 414804 596476 415404 596478
rect 450804 596476 451404 596478
rect 486804 596476 487404 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586260 596476 586860 596478
rect -2936 596454 586860 596476
rect -2936 596218 -2754 596454
rect -2518 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 90986 596454
rect 91222 596218 126986 596454
rect 127222 596218 162986 596454
rect 163222 596218 198986 596454
rect 199222 596218 234986 596454
rect 235222 596218 270986 596454
rect 271222 596218 306986 596454
rect 307222 596218 342986 596454
rect 343222 596218 378986 596454
rect 379222 596218 414986 596454
rect 415222 596218 450986 596454
rect 451222 596218 486986 596454
rect 487222 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586442 596454
rect 586678 596218 586860 596454
rect -2936 596134 586860 596218
rect -2936 595898 -2754 596134
rect -2518 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 90986 596134
rect 91222 595898 126986 596134
rect 127222 595898 162986 596134
rect 163222 595898 198986 596134
rect 199222 595898 234986 596134
rect 235222 595898 270986 596134
rect 271222 595898 306986 596134
rect 307222 595898 342986 596134
rect 343222 595898 378986 596134
rect 379222 595898 414986 596134
rect 415222 595898 450986 596134
rect 451222 595898 486986 596134
rect 487222 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586442 596134
rect 586678 595898 586860 596134
rect -2936 595876 586860 595898
rect -2936 595874 -2336 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 90804 595874 91404 595876
rect 126804 595874 127404 595876
rect 162804 595874 163404 595876
rect 198804 595874 199404 595876
rect 234804 595874 235404 595876
rect 270804 595874 271404 595876
rect 306804 595874 307404 595876
rect 342804 595874 343404 595876
rect 378804 595874 379404 595876
rect 414804 595874 415404 595876
rect 450804 595874 451404 595876
rect 486804 595874 487404 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586260 595874 586860 595876
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 262128 578476 262448 578478
rect 288804 578476 289404 578478
rect 554256 578476 554576 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2936 578454 586860 578476
rect -2936 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 262170 578454
rect 262406 578218 288986 578454
rect 289222 578218 554298 578454
rect 554534 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586860 578454
rect -2936 578134 586860 578218
rect -2936 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 262170 578134
rect 262406 577898 288986 578134
rect 289222 577898 554298 578134
rect 554534 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586860 578134
rect -2936 577876 586860 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 262128 577874 262448 577876
rect 288804 577874 289404 577876
rect 554256 577874 554576 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -2936 560476 -2336 560478
rect 18804 560476 19404 560478
rect 246768 560476 247088 560478
rect 270804 560476 271404 560478
rect 306804 560476 307404 560478
rect 538896 560476 539216 560478
rect 586260 560476 586860 560478
rect -2936 560454 586860 560476
rect -2936 560218 -2754 560454
rect -2518 560218 18986 560454
rect 19222 560218 246810 560454
rect 247046 560218 270986 560454
rect 271222 560218 306986 560454
rect 307222 560218 538938 560454
rect 539174 560218 586442 560454
rect 586678 560218 586860 560454
rect -2936 560134 586860 560218
rect -2936 559898 -2754 560134
rect -2518 559898 18986 560134
rect 19222 559898 246810 560134
rect 247046 559898 270986 560134
rect 271222 559898 306986 560134
rect 307222 559898 538938 560134
rect 539174 559898 586442 560134
rect 586678 559898 586860 560134
rect -2936 559876 586860 559898
rect -2936 559874 -2336 559876
rect 18804 559874 19404 559876
rect 246768 559874 247088 559876
rect 270804 559874 271404 559876
rect 306804 559874 307404 559876
rect 538896 559874 539216 559876
rect 586260 559874 586860 559876
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 262128 542476 262448 542478
rect 288804 542476 289404 542478
rect 554256 542476 554576 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2936 542454 586860 542476
rect -2936 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 262170 542454
rect 262406 542218 288986 542454
rect 289222 542218 554298 542454
rect 554534 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586860 542454
rect -2936 542134 586860 542218
rect -2936 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 262170 542134
rect 262406 541898 288986 542134
rect 289222 541898 554298 542134
rect 554534 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586860 542134
rect -2936 541876 586860 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 262128 541874 262448 541876
rect 288804 541874 289404 541876
rect 554256 541874 554576 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -2936 524476 -2336 524478
rect 18804 524476 19404 524478
rect 246768 524476 247088 524478
rect 270804 524476 271404 524478
rect 306804 524476 307404 524478
rect 538896 524476 539216 524478
rect 586260 524476 586860 524478
rect -2936 524454 586860 524476
rect -2936 524218 -2754 524454
rect -2518 524218 18986 524454
rect 19222 524218 246810 524454
rect 247046 524218 270986 524454
rect 271222 524218 306986 524454
rect 307222 524218 538938 524454
rect 539174 524218 586442 524454
rect 586678 524218 586860 524454
rect -2936 524134 586860 524218
rect -2936 523898 -2754 524134
rect -2518 523898 18986 524134
rect 19222 523898 246810 524134
rect 247046 523898 270986 524134
rect 271222 523898 306986 524134
rect 307222 523898 538938 524134
rect 539174 523898 586442 524134
rect 586678 523898 586860 524134
rect -2936 523876 586860 523898
rect -2936 523874 -2336 523876
rect 18804 523874 19404 523876
rect 246768 523874 247088 523876
rect 270804 523874 271404 523876
rect 306804 523874 307404 523876
rect 538896 523874 539216 523876
rect 586260 523874 586860 523876
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 262128 506476 262448 506478
rect 288804 506476 289404 506478
rect 554256 506476 554576 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2936 506454 586860 506476
rect -2936 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 262170 506454
rect 262406 506218 288986 506454
rect 289222 506218 554298 506454
rect 554534 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586860 506454
rect -2936 506134 586860 506218
rect -2936 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 262170 506134
rect 262406 505898 288986 506134
rect 289222 505898 554298 506134
rect 554534 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586860 506134
rect -2936 505876 586860 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 262128 505874 262448 505876
rect 288804 505874 289404 505876
rect 554256 505874 554576 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -2936 488476 -2336 488478
rect 18804 488476 19404 488478
rect 246768 488476 247088 488478
rect 270804 488476 271404 488478
rect 306804 488476 307404 488478
rect 538896 488476 539216 488478
rect 586260 488476 586860 488478
rect -2936 488454 586860 488476
rect -2936 488218 -2754 488454
rect -2518 488218 18986 488454
rect 19222 488218 246810 488454
rect 247046 488218 270986 488454
rect 271222 488218 306986 488454
rect 307222 488218 538938 488454
rect 539174 488218 586442 488454
rect 586678 488218 586860 488454
rect -2936 488134 586860 488218
rect -2936 487898 -2754 488134
rect -2518 487898 18986 488134
rect 19222 487898 246810 488134
rect 247046 487898 270986 488134
rect 271222 487898 306986 488134
rect 307222 487898 538938 488134
rect 539174 487898 586442 488134
rect 586678 487898 586860 488134
rect -2936 487876 586860 487898
rect -2936 487874 -2336 487876
rect 18804 487874 19404 487876
rect 246768 487874 247088 487876
rect 270804 487874 271404 487876
rect 306804 487874 307404 487876
rect 538896 487874 539216 487876
rect 586260 487874 586860 487876
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 262128 470476 262448 470478
rect 288804 470476 289404 470478
rect 554256 470476 554576 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2936 470454 586860 470476
rect -2936 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 262170 470454
rect 262406 470218 288986 470454
rect 289222 470218 554298 470454
rect 554534 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586860 470454
rect -2936 470134 586860 470218
rect -2936 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 262170 470134
rect 262406 469898 288986 470134
rect 289222 469898 554298 470134
rect 554534 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586860 470134
rect -2936 469876 586860 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 262128 469874 262448 469876
rect 288804 469874 289404 469876
rect 554256 469874 554576 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -2936 452476 -2336 452478
rect 18804 452476 19404 452478
rect 246768 452476 247088 452478
rect 270804 452476 271404 452478
rect 306804 452476 307404 452478
rect 538896 452476 539216 452478
rect 586260 452476 586860 452478
rect -2936 452454 586860 452476
rect -2936 452218 -2754 452454
rect -2518 452218 18986 452454
rect 19222 452218 246810 452454
rect 247046 452218 270986 452454
rect 271222 452218 306986 452454
rect 307222 452218 538938 452454
rect 539174 452218 586442 452454
rect 586678 452218 586860 452454
rect -2936 452134 586860 452218
rect -2936 451898 -2754 452134
rect -2518 451898 18986 452134
rect 19222 451898 246810 452134
rect 247046 451898 270986 452134
rect 271222 451898 306986 452134
rect 307222 451898 538938 452134
rect 539174 451898 586442 452134
rect 586678 451898 586860 452134
rect -2936 451876 586860 451898
rect -2936 451874 -2336 451876
rect 18804 451874 19404 451876
rect 246768 451874 247088 451876
rect 270804 451874 271404 451876
rect 306804 451874 307404 451876
rect 538896 451874 539216 451876
rect 586260 451874 586860 451876
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 262128 434476 262448 434478
rect 288804 434476 289404 434478
rect 554256 434476 554576 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2936 434454 586860 434476
rect -2936 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 262170 434454
rect 262406 434218 288986 434454
rect 289222 434218 554298 434454
rect 554534 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586860 434454
rect -2936 434134 586860 434218
rect -2936 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 262170 434134
rect 262406 433898 288986 434134
rect 289222 433898 554298 434134
rect 554534 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586860 434134
rect -2936 433876 586860 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 262128 433874 262448 433876
rect 288804 433874 289404 433876
rect 554256 433874 554576 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -2936 416476 -2336 416478
rect 18804 416476 19404 416478
rect 246768 416476 247088 416478
rect 270804 416476 271404 416478
rect 306804 416476 307404 416478
rect 538896 416476 539216 416478
rect 586260 416476 586860 416478
rect -2936 416454 586860 416476
rect -2936 416218 -2754 416454
rect -2518 416218 18986 416454
rect 19222 416218 246810 416454
rect 247046 416218 270986 416454
rect 271222 416218 306986 416454
rect 307222 416218 538938 416454
rect 539174 416218 586442 416454
rect 586678 416218 586860 416454
rect -2936 416134 586860 416218
rect -2936 415898 -2754 416134
rect -2518 415898 18986 416134
rect 19222 415898 246810 416134
rect 247046 415898 270986 416134
rect 271222 415898 306986 416134
rect 307222 415898 538938 416134
rect 539174 415898 586442 416134
rect 586678 415898 586860 416134
rect -2936 415876 586860 415898
rect -2936 415874 -2336 415876
rect 18804 415874 19404 415876
rect 246768 415874 247088 415876
rect 270804 415874 271404 415876
rect 306804 415874 307404 415876
rect 538896 415874 539216 415876
rect 586260 415874 586860 415876
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 262128 398476 262448 398478
rect 288804 398476 289404 398478
rect 554256 398476 554576 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2936 398454 586860 398476
rect -2936 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 262170 398454
rect 262406 398218 288986 398454
rect 289222 398218 554298 398454
rect 554534 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586860 398454
rect -2936 398134 586860 398218
rect -2936 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 262170 398134
rect 262406 397898 288986 398134
rect 289222 397898 554298 398134
rect 554534 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586860 398134
rect -2936 397876 586860 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 262128 397874 262448 397876
rect 288804 397874 289404 397876
rect 554256 397874 554576 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -2936 380476 -2336 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 90804 380476 91404 380478
rect 126804 380476 127404 380478
rect 162804 380476 163404 380478
rect 198804 380476 199404 380478
rect 234804 380476 235404 380478
rect 270804 380476 271404 380478
rect 306804 380476 307404 380478
rect 342804 380476 343404 380478
rect 378804 380476 379404 380478
rect 414804 380476 415404 380478
rect 450804 380476 451404 380478
rect 486804 380476 487404 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586260 380476 586860 380478
rect -2936 380454 586860 380476
rect -2936 380218 -2754 380454
rect -2518 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 90986 380454
rect 91222 380218 126986 380454
rect 127222 380218 162986 380454
rect 163222 380218 198986 380454
rect 199222 380218 234986 380454
rect 235222 380218 270986 380454
rect 271222 380218 306986 380454
rect 307222 380218 342986 380454
rect 343222 380218 378986 380454
rect 379222 380218 414986 380454
rect 415222 380218 450986 380454
rect 451222 380218 486986 380454
rect 487222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586442 380454
rect 586678 380218 586860 380454
rect -2936 380134 586860 380218
rect -2936 379898 -2754 380134
rect -2518 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 90986 380134
rect 91222 379898 126986 380134
rect 127222 379898 162986 380134
rect 163222 379898 198986 380134
rect 199222 379898 234986 380134
rect 235222 379898 270986 380134
rect 271222 379898 306986 380134
rect 307222 379898 342986 380134
rect 343222 379898 378986 380134
rect 379222 379898 414986 380134
rect 415222 379898 450986 380134
rect 451222 379898 486986 380134
rect 487222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586442 380134
rect 586678 379898 586860 380134
rect -2936 379876 586860 379898
rect -2936 379874 -2336 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 90804 379874 91404 379876
rect 126804 379874 127404 379876
rect 162804 379874 163404 379876
rect 198804 379874 199404 379876
rect 234804 379874 235404 379876
rect 270804 379874 271404 379876
rect 306804 379874 307404 379876
rect 342804 379874 343404 379876
rect 378804 379874 379404 379876
rect 414804 379874 415404 379876
rect 450804 379874 451404 379876
rect 486804 379874 487404 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586260 379874 586860 379876
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 72804 362476 73404 362478
rect 108804 362476 109404 362478
rect 144804 362476 145404 362478
rect 180804 362476 181404 362478
rect 216804 362476 217404 362478
rect 252804 362476 253404 362478
rect 288804 362476 289404 362478
rect 324804 362476 325404 362478
rect 360804 362476 361404 362478
rect 396804 362476 397404 362478
rect 432804 362476 433404 362478
rect 468804 362476 469404 362478
rect 504804 362476 505404 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2936 362454 586860 362476
rect -2936 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 72986 362454
rect 73222 362218 108986 362454
rect 109222 362218 144986 362454
rect 145222 362218 180986 362454
rect 181222 362218 216986 362454
rect 217222 362218 252986 362454
rect 253222 362218 288986 362454
rect 289222 362218 324986 362454
rect 325222 362218 360986 362454
rect 361222 362218 396986 362454
rect 397222 362218 432986 362454
rect 433222 362218 468986 362454
rect 469222 362218 504986 362454
rect 505222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586860 362454
rect -2936 362134 586860 362218
rect -2936 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 72986 362134
rect 73222 361898 108986 362134
rect 109222 361898 144986 362134
rect 145222 361898 180986 362134
rect 181222 361898 216986 362134
rect 217222 361898 252986 362134
rect 253222 361898 288986 362134
rect 289222 361898 324986 362134
rect 325222 361898 360986 362134
rect 361222 361898 396986 362134
rect 397222 361898 432986 362134
rect 433222 361898 468986 362134
rect 469222 361898 504986 362134
rect 505222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586860 362134
rect -2936 361876 586860 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 72804 361874 73404 361876
rect 108804 361874 109404 361876
rect 144804 361874 145404 361876
rect 180804 361874 181404 361876
rect 216804 361874 217404 361876
rect 252804 361874 253404 361876
rect 288804 361874 289404 361876
rect 324804 361874 325404 361876
rect 360804 361874 361404 361876
rect 396804 361874 397404 361876
rect 432804 361874 433404 361876
rect 468804 361874 469404 361876
rect 504804 361874 505404 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -2936 344476 -2336 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 90804 344476 91404 344478
rect 126804 344476 127404 344478
rect 162804 344476 163404 344478
rect 198804 344476 199404 344478
rect 234804 344476 235404 344478
rect 292112 344476 292432 344478
rect 342804 344476 343404 344478
rect 378804 344476 379404 344478
rect 414804 344476 415404 344478
rect 450804 344476 451404 344478
rect 486804 344476 487404 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586260 344476 586860 344478
rect -2936 344454 586860 344476
rect -2936 344218 -2754 344454
rect -2518 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 90986 344454
rect 91222 344218 126986 344454
rect 127222 344218 162986 344454
rect 163222 344218 198986 344454
rect 199222 344218 234986 344454
rect 235222 344218 292154 344454
rect 292390 344218 342986 344454
rect 343222 344218 378986 344454
rect 379222 344218 414986 344454
rect 415222 344218 450986 344454
rect 451222 344218 486986 344454
rect 487222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586442 344454
rect 586678 344218 586860 344454
rect -2936 344134 586860 344218
rect -2936 343898 -2754 344134
rect -2518 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 90986 344134
rect 91222 343898 126986 344134
rect 127222 343898 162986 344134
rect 163222 343898 198986 344134
rect 199222 343898 234986 344134
rect 235222 343898 292154 344134
rect 292390 343898 342986 344134
rect 343222 343898 378986 344134
rect 379222 343898 414986 344134
rect 415222 343898 450986 344134
rect 451222 343898 486986 344134
rect 487222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586442 344134
rect 586678 343898 586860 344134
rect -2936 343876 586860 343898
rect -2936 343874 -2336 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 90804 343874 91404 343876
rect 126804 343874 127404 343876
rect 162804 343874 163404 343876
rect 198804 343874 199404 343876
rect 234804 343874 235404 343876
rect 292112 343874 292432 343876
rect 342804 343874 343404 343876
rect 378804 343874 379404 343876
rect 414804 343874 415404 343876
rect 450804 343874 451404 343876
rect 486804 343874 487404 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586260 343874 586860 343876
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 72804 326476 73404 326478
rect 108804 326476 109404 326478
rect 144804 326476 145404 326478
rect 180804 326476 181404 326478
rect 216804 326476 217404 326478
rect 252804 326476 253404 326478
rect 307472 326476 307792 326478
rect 324804 326476 325404 326478
rect 360804 326476 361404 326478
rect 396804 326476 397404 326478
rect 432804 326476 433404 326478
rect 468804 326476 469404 326478
rect 504804 326476 505404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2936 326454 586860 326476
rect -2936 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 72986 326454
rect 73222 326218 108986 326454
rect 109222 326218 144986 326454
rect 145222 326218 180986 326454
rect 181222 326218 216986 326454
rect 217222 326218 252986 326454
rect 253222 326218 307514 326454
rect 307750 326218 324986 326454
rect 325222 326218 360986 326454
rect 361222 326218 396986 326454
rect 397222 326218 432986 326454
rect 433222 326218 468986 326454
rect 469222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586860 326454
rect -2936 326134 586860 326218
rect -2936 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 72986 326134
rect 73222 325898 108986 326134
rect 109222 325898 144986 326134
rect 145222 325898 180986 326134
rect 181222 325898 216986 326134
rect 217222 325898 252986 326134
rect 253222 325898 307514 326134
rect 307750 325898 324986 326134
rect 325222 325898 360986 326134
rect 361222 325898 396986 326134
rect 397222 325898 432986 326134
rect 433222 325898 468986 326134
rect 469222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586860 326134
rect -2936 325876 586860 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 72804 325874 73404 325876
rect 108804 325874 109404 325876
rect 144804 325874 145404 325876
rect 180804 325874 181404 325876
rect 216804 325874 217404 325876
rect 252804 325874 253404 325876
rect 307472 325874 307792 325876
rect 324804 325874 325404 325876
rect 360804 325874 361404 325876
rect 396804 325874 397404 325876
rect 432804 325874 433404 325876
rect 468804 325874 469404 325876
rect 504804 325874 505404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -2936 308476 -2336 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 90804 308476 91404 308478
rect 126804 308476 127404 308478
rect 162804 308476 163404 308478
rect 198804 308476 199404 308478
rect 234804 308476 235404 308478
rect 270804 308476 271404 308478
rect 306804 308476 307404 308478
rect 342804 308476 343404 308478
rect 378804 308476 379404 308478
rect 414804 308476 415404 308478
rect 450804 308476 451404 308478
rect 486804 308476 487404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586260 308476 586860 308478
rect -2936 308454 586860 308476
rect -2936 308218 -2754 308454
rect -2518 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 90986 308454
rect 91222 308218 126986 308454
rect 127222 308218 162986 308454
rect 163222 308218 198986 308454
rect 199222 308218 234986 308454
rect 235222 308218 270986 308454
rect 271222 308218 306986 308454
rect 307222 308218 342986 308454
rect 343222 308218 378986 308454
rect 379222 308218 414986 308454
rect 415222 308218 450986 308454
rect 451222 308218 486986 308454
rect 487222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586442 308454
rect 586678 308218 586860 308454
rect -2936 308134 586860 308218
rect -2936 307898 -2754 308134
rect -2518 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 90986 308134
rect 91222 307898 126986 308134
rect 127222 307898 162986 308134
rect 163222 307898 198986 308134
rect 199222 307898 234986 308134
rect 235222 307898 270986 308134
rect 271222 307898 306986 308134
rect 307222 307898 342986 308134
rect 343222 307898 378986 308134
rect 379222 307898 414986 308134
rect 415222 307898 450986 308134
rect 451222 307898 486986 308134
rect 487222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586442 308134
rect 586678 307898 586860 308134
rect -2936 307876 586860 307898
rect -2936 307874 -2336 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 90804 307874 91404 307876
rect 126804 307874 127404 307876
rect 162804 307874 163404 307876
rect 198804 307874 199404 307876
rect 234804 307874 235404 307876
rect 270804 307874 271404 307876
rect 306804 307874 307404 307876
rect 342804 307874 343404 307876
rect 378804 307874 379404 307876
rect 414804 307874 415404 307876
rect 450804 307874 451404 307876
rect 486804 307874 487404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586260 307874 586860 307876
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 108804 290476 109404 290478
rect 144804 290476 145404 290478
rect 180804 290476 181404 290478
rect 216804 290476 217404 290478
rect 252804 290476 253404 290478
rect 288804 290476 289404 290478
rect 324804 290476 325404 290478
rect 360804 290476 361404 290478
rect 396804 290476 397404 290478
rect 432804 290476 433404 290478
rect 468804 290476 469404 290478
rect 504804 290476 505404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2936 290454 586860 290476
rect -2936 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 108986 290454
rect 109222 290218 144986 290454
rect 145222 290218 180986 290454
rect 181222 290218 216986 290454
rect 217222 290218 252986 290454
rect 253222 290218 288986 290454
rect 289222 290218 324986 290454
rect 325222 290218 360986 290454
rect 361222 290218 396986 290454
rect 397222 290218 432986 290454
rect 433222 290218 468986 290454
rect 469222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586860 290454
rect -2936 290134 586860 290218
rect -2936 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 108986 290134
rect 109222 289898 144986 290134
rect 145222 289898 180986 290134
rect 181222 289898 216986 290134
rect 217222 289898 252986 290134
rect 253222 289898 288986 290134
rect 289222 289898 324986 290134
rect 325222 289898 360986 290134
rect 361222 289898 396986 290134
rect 397222 289898 432986 290134
rect 433222 289898 468986 290134
rect 469222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586860 290134
rect -2936 289876 586860 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 108804 289874 109404 289876
rect 144804 289874 145404 289876
rect 180804 289874 181404 289876
rect 216804 289874 217404 289876
rect 252804 289874 253404 289876
rect 288804 289874 289404 289876
rect 324804 289874 325404 289876
rect 360804 289874 361404 289876
rect 396804 289874 397404 289876
rect 432804 289874 433404 289876
rect 468804 289874 469404 289876
rect 504804 289874 505404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -2936 272476 -2336 272478
rect 18804 272476 19404 272478
rect 270804 272476 271404 272478
rect 306804 272476 307404 272478
rect 586260 272476 586860 272478
rect -2936 272454 586860 272476
rect -2936 272218 -2754 272454
rect -2518 272218 18986 272454
rect 19222 272218 270986 272454
rect 271222 272218 306986 272454
rect 307222 272218 586442 272454
rect 586678 272218 586860 272454
rect -2936 272134 586860 272218
rect -2936 271898 -2754 272134
rect -2518 271898 18986 272134
rect 19222 271898 270986 272134
rect 271222 271898 306986 272134
rect 307222 271898 586442 272134
rect 586678 271898 586860 272134
rect -2936 271876 586860 271898
rect -2936 271874 -2336 271876
rect 18804 271874 19404 271876
rect 270804 271874 271404 271876
rect 306804 271874 307404 271876
rect 586260 271874 586860 271876
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 262128 254476 262448 254478
rect 288804 254476 289404 254478
rect 554256 254476 554576 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2936 254454 586860 254476
rect -2936 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 262170 254454
rect 262406 254218 288986 254454
rect 289222 254218 554298 254454
rect 554534 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586860 254454
rect -2936 254134 586860 254218
rect -2936 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 262170 254134
rect 262406 253898 288986 254134
rect 289222 253898 554298 254134
rect 554534 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586860 254134
rect -2936 253876 586860 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 262128 253874 262448 253876
rect 288804 253874 289404 253876
rect 554256 253874 554576 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -2936 236476 -2336 236478
rect 18804 236476 19404 236478
rect 246768 236476 247088 236478
rect 270804 236476 271404 236478
rect 306804 236476 307404 236478
rect 538896 236476 539216 236478
rect 586260 236476 586860 236478
rect -2936 236454 586860 236476
rect -2936 236218 -2754 236454
rect -2518 236218 18986 236454
rect 19222 236218 246810 236454
rect 247046 236218 270986 236454
rect 271222 236218 306986 236454
rect 307222 236218 538938 236454
rect 539174 236218 586442 236454
rect 586678 236218 586860 236454
rect -2936 236134 586860 236218
rect -2936 235898 -2754 236134
rect -2518 235898 18986 236134
rect 19222 235898 246810 236134
rect 247046 235898 270986 236134
rect 271222 235898 306986 236134
rect 307222 235898 538938 236134
rect 539174 235898 586442 236134
rect 586678 235898 586860 236134
rect -2936 235876 586860 235898
rect -2936 235874 -2336 235876
rect 18804 235874 19404 235876
rect 246768 235874 247088 235876
rect 270804 235874 271404 235876
rect 306804 235874 307404 235876
rect 538896 235874 539216 235876
rect 586260 235874 586860 235876
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 262128 218476 262448 218478
rect 288804 218476 289404 218478
rect 554256 218476 554576 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2936 218454 586860 218476
rect -2936 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 262170 218454
rect 262406 218218 288986 218454
rect 289222 218218 554298 218454
rect 554534 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586860 218454
rect -2936 218134 586860 218218
rect -2936 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 262170 218134
rect 262406 217898 288986 218134
rect 289222 217898 554298 218134
rect 554534 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586860 218134
rect -2936 217876 586860 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 262128 217874 262448 217876
rect 288804 217874 289404 217876
rect 554256 217874 554576 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -2936 200476 -2336 200478
rect 18804 200476 19404 200478
rect 246768 200476 247088 200478
rect 270804 200476 271404 200478
rect 306804 200476 307404 200478
rect 538896 200476 539216 200478
rect 586260 200476 586860 200478
rect -2936 200454 586860 200476
rect -2936 200218 -2754 200454
rect -2518 200218 18986 200454
rect 19222 200218 246810 200454
rect 247046 200218 270986 200454
rect 271222 200218 306986 200454
rect 307222 200218 538938 200454
rect 539174 200218 586442 200454
rect 586678 200218 586860 200454
rect -2936 200134 586860 200218
rect -2936 199898 -2754 200134
rect -2518 199898 18986 200134
rect 19222 199898 246810 200134
rect 247046 199898 270986 200134
rect 271222 199898 306986 200134
rect 307222 199898 538938 200134
rect 539174 199898 586442 200134
rect 586678 199898 586860 200134
rect -2936 199876 586860 199898
rect -2936 199874 -2336 199876
rect 18804 199874 19404 199876
rect 246768 199874 247088 199876
rect 270804 199874 271404 199876
rect 306804 199874 307404 199876
rect 538896 199874 539216 199876
rect 586260 199874 586860 199876
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 262128 182476 262448 182478
rect 288804 182476 289404 182478
rect 554256 182476 554576 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2936 182454 586860 182476
rect -2936 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 262170 182454
rect 262406 182218 288986 182454
rect 289222 182218 554298 182454
rect 554534 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586860 182454
rect -2936 182134 586860 182218
rect -2936 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 262170 182134
rect 262406 181898 288986 182134
rect 289222 181898 554298 182134
rect 554534 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586860 182134
rect -2936 181876 586860 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 262128 181874 262448 181876
rect 288804 181874 289404 181876
rect 554256 181874 554576 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -2936 164476 -2336 164478
rect 18804 164476 19404 164478
rect 246768 164476 247088 164478
rect 270804 164476 271404 164478
rect 306804 164476 307404 164478
rect 538896 164476 539216 164478
rect 586260 164476 586860 164478
rect -2936 164454 586860 164476
rect -2936 164218 -2754 164454
rect -2518 164218 18986 164454
rect 19222 164218 246810 164454
rect 247046 164218 270986 164454
rect 271222 164218 306986 164454
rect 307222 164218 538938 164454
rect 539174 164218 586442 164454
rect 586678 164218 586860 164454
rect -2936 164134 586860 164218
rect -2936 163898 -2754 164134
rect -2518 163898 18986 164134
rect 19222 163898 246810 164134
rect 247046 163898 270986 164134
rect 271222 163898 306986 164134
rect 307222 163898 538938 164134
rect 539174 163898 586442 164134
rect 586678 163898 586860 164134
rect -2936 163876 586860 163898
rect -2936 163874 -2336 163876
rect 18804 163874 19404 163876
rect 246768 163874 247088 163876
rect 270804 163874 271404 163876
rect 306804 163874 307404 163876
rect 538896 163874 539216 163876
rect 586260 163874 586860 163876
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 262128 146476 262448 146478
rect 288804 146476 289404 146478
rect 554256 146476 554576 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2936 146454 586860 146476
rect -2936 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 262170 146454
rect 262406 146218 288986 146454
rect 289222 146218 554298 146454
rect 554534 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586860 146454
rect -2936 146134 586860 146218
rect -2936 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 262170 146134
rect 262406 145898 288986 146134
rect 289222 145898 554298 146134
rect 554534 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586860 146134
rect -2936 145876 586860 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 262128 145874 262448 145876
rect 288804 145874 289404 145876
rect 554256 145874 554576 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -2936 128476 -2336 128478
rect 18804 128476 19404 128478
rect 246768 128476 247088 128478
rect 270804 128476 271404 128478
rect 306804 128476 307404 128478
rect 538896 128476 539216 128478
rect 586260 128476 586860 128478
rect -2936 128454 586860 128476
rect -2936 128218 -2754 128454
rect -2518 128218 18986 128454
rect 19222 128218 246810 128454
rect 247046 128218 270986 128454
rect 271222 128218 306986 128454
rect 307222 128218 538938 128454
rect 539174 128218 586442 128454
rect 586678 128218 586860 128454
rect -2936 128134 586860 128218
rect -2936 127898 -2754 128134
rect -2518 127898 18986 128134
rect 19222 127898 246810 128134
rect 247046 127898 270986 128134
rect 271222 127898 306986 128134
rect 307222 127898 538938 128134
rect 539174 127898 586442 128134
rect 586678 127898 586860 128134
rect -2936 127876 586860 127898
rect -2936 127874 -2336 127876
rect 18804 127874 19404 127876
rect 246768 127874 247088 127876
rect 270804 127874 271404 127876
rect 306804 127874 307404 127876
rect 538896 127874 539216 127876
rect 586260 127874 586860 127876
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 262128 110476 262448 110478
rect 288804 110476 289404 110478
rect 554256 110476 554576 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2936 110454 586860 110476
rect -2936 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 262170 110454
rect 262406 110218 288986 110454
rect 289222 110218 554298 110454
rect 554534 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586860 110454
rect -2936 110134 586860 110218
rect -2936 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 262170 110134
rect 262406 109898 288986 110134
rect 289222 109898 554298 110134
rect 554534 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586860 110134
rect -2936 109876 586860 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 262128 109874 262448 109876
rect 288804 109874 289404 109876
rect 554256 109874 554576 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -2936 92476 -2336 92478
rect 18804 92476 19404 92478
rect 246768 92476 247088 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 538896 92476 539216 92478
rect 586260 92476 586860 92478
rect -2936 92454 586860 92476
rect -2936 92218 -2754 92454
rect -2518 92218 18986 92454
rect 19222 92218 246810 92454
rect 247046 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 538938 92454
rect 539174 92218 586442 92454
rect 586678 92218 586860 92454
rect -2936 92134 586860 92218
rect -2936 91898 -2754 92134
rect -2518 91898 18986 92134
rect 19222 91898 246810 92134
rect 247046 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 538938 92134
rect 539174 91898 586442 92134
rect 586678 91898 586860 92134
rect -2936 91876 586860 91898
rect -2936 91874 -2336 91876
rect 18804 91874 19404 91876
rect 246768 91874 247088 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 538896 91874 539216 91876
rect 586260 91874 586860 91876
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 288804 74476 289404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2936 74454 586860 74476
rect -2936 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 288986 74454
rect 289222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586860 74454
rect -2936 74134 586860 74218
rect -2936 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 288986 74134
rect 289222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586860 74134
rect -2936 73876 586860 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 288804 73874 289404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -2936 56476 -2336 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586260 56476 586860 56478
rect -2936 56454 586860 56476
rect -2936 56218 -2754 56454
rect -2518 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586442 56454
rect 586678 56218 586860 56454
rect -2936 56134 586860 56218
rect -2936 55898 -2754 56134
rect -2518 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586442 56134
rect 586678 55898 586860 56134
rect -2936 55876 586860 55898
rect -2936 55874 -2336 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586260 55874 586860 55876
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2936 38454 586860 38476
rect -2936 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586860 38454
rect -2936 38134 586860 38218
rect -2936 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586860 38134
rect -2936 37876 586860 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -2936 20476 -2336 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586260 20476 586860 20478
rect -2936 20454 586860 20476
rect -2936 20218 -2754 20454
rect -2518 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586442 20454
rect 586678 20218 586860 20454
rect -2936 20134 586860 20218
rect -2936 19898 -2754 20134
rect -2518 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586442 20134
rect 586678 19898 586860 20134
rect -2936 19876 586860 19898
rect -2936 19874 -2336 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586260 19874 586860 19876
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2936 2454 586860 2476
rect -2936 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586860 2454
rect -2936 2134 586860 2218
rect -2936 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586860 2134
rect -2936 1876 586860 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 18804 -1264 19404 -1262
rect 54804 -1264 55404 -1262
rect 90804 -1264 91404 -1262
rect 126804 -1264 127404 -1262
rect 162804 -1264 163404 -1262
rect 198804 -1264 199404 -1262
rect 234804 -1264 235404 -1262
rect 270804 -1264 271404 -1262
rect 306804 -1264 307404 -1262
rect 342804 -1264 343404 -1262
rect 378804 -1264 379404 -1262
rect 414804 -1264 415404 -1262
rect 450804 -1264 451404 -1262
rect 486804 -1264 487404 -1262
rect 522804 -1264 523404 -1262
rect 558804 -1264 559404 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1286 586860 -1264
rect -2936 -1522 -2754 -1286
rect -2518 -1522 18986 -1286
rect 19222 -1522 54986 -1286
rect 55222 -1522 90986 -1286
rect 91222 -1522 126986 -1286
rect 127222 -1522 162986 -1286
rect 163222 -1522 198986 -1286
rect 199222 -1522 234986 -1286
rect 235222 -1522 270986 -1286
rect 271222 -1522 306986 -1286
rect 307222 -1522 342986 -1286
rect 343222 -1522 378986 -1286
rect 379222 -1522 414986 -1286
rect 415222 -1522 450986 -1286
rect 451222 -1522 486986 -1286
rect 487222 -1522 522986 -1286
rect 523222 -1522 558986 -1286
rect 559222 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect -2936 -1606 586860 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 18986 -1606
rect 19222 -1842 54986 -1606
rect 55222 -1842 90986 -1606
rect 91222 -1842 126986 -1606
rect 127222 -1842 162986 -1606
rect 163222 -1842 198986 -1606
rect 199222 -1842 234986 -1606
rect 235222 -1842 270986 -1606
rect 271222 -1842 306986 -1606
rect 307222 -1842 342986 -1606
rect 343222 -1842 378986 -1606
rect 379222 -1842 414986 -1606
rect 415222 -1842 450986 -1606
rect 451222 -1842 486986 -1606
rect 487222 -1842 522986 -1606
rect 523222 -1842 558986 -1606
rect 559222 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect -2936 -1864 586860 -1842
rect -2936 -1866 -2336 -1864
rect 18804 -1866 19404 -1864
rect 54804 -1866 55404 -1864
rect 90804 -1866 91404 -1864
rect 126804 -1866 127404 -1864
rect 162804 -1866 163404 -1864
rect 198804 -1866 199404 -1864
rect 234804 -1866 235404 -1864
rect 270804 -1866 271404 -1864
rect 306804 -1866 307404 -1864
rect 342804 -1866 343404 -1864
rect 378804 -1866 379404 -1864
rect 414804 -1866 415404 -1864
rect 450804 -1866 451404 -1864
rect 486804 -1866 487404 -1864
rect 522804 -1866 523404 -1864
rect 558804 -1866 559404 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2226 587800 -2204
rect -3876 -2462 -3694 -2226
rect -3458 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect -3876 -2546 587800 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect -3876 -2804 587800 -2782
rect -3876 -2806 -3276 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3166 588740 -3144
rect -4816 -3402 -4634 -3166
rect -4398 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect -4816 -3486 588740 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect -4816 -3744 588740 -3722
rect -4816 -3746 -4216 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4106 589680 -4084
rect -5756 -4342 -5574 -4106
rect -5338 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect -5756 -4426 589680 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect -5756 -4684 589680 -4662
rect -5756 -4686 -5156 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5046 590620 -5024
rect -6696 -5282 -6514 -5046
rect -6278 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect -6696 -5366 590620 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect -6696 -5624 590620 -5602
rect -6696 -5626 -6096 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 590960 -5964 591560 -5962
rect -7636 -5986 591560 -5964
rect -7636 -6222 -7454 -5986
rect -7218 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect -7636 -6306 591560 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect -7636 -6564 591560 -6542
rect -7636 -6566 -7036 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 591900 -6904 592500 -6902
rect -8576 -6926 592500 -6904
rect -8576 -7162 -8394 -6926
rect -8158 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect -8576 -7246 592500 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect -8576 -7504 592500 -7482
rect -8576 -7506 -7976 -7504
rect 591900 -7506 592500 -7504
use decred_hash_macro  decred_hash_block3
timestamp 1608091038
transform -1 0 558784 0 -1 583916
box 0 0 240000 200000
use decred_hash_macro  decred_hash_block2
timestamp 1608091038
transform -1 0 266656 0 -1 583916
box 0 0 240000 200000
use decred_hash_macro  decred_hash_block1
timestamp 1608091038
transform -1 0 558784 0 -1 273600
box 0 0 240000 200000
use decred_hash_macro  decred_hash_block0
timestamp 1608091038
transform -1 0 266656 0 -1 273600
box 0 0 240000 200000
use decred_controller  decred_controller_block
timestamp 1608091038
transform -1 0 312000 0 -1 355560
box 0 0 40000 40000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 70 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 71 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 72 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 73 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 74 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 75 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 76 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 77 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 78 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 79 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 80 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 81 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 82 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 83 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 84 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 85 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 86 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 87 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 88 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 89 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 90 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 91 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 92 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 93 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 94 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 95 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 96 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 97 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 98 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 99 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 100 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 101 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 102 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 103 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 104 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 105 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 106 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 107 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 108 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 109 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 110 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 111 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 112 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 113 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 114 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 115 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 116 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 117 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 118 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 119 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 120 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 121 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 122 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 123 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 124 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 125 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 126 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 127 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 128 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 129 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 130 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 131 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 132 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 133 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 134 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 135 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 136 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 137 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 138 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 139 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 140 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 141 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 142 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 143 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 144 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 145 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 146 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 147 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 148 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 149 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 150 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 151 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 152 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 153 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 154 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 155 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 156 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 157 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 158 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 159 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 160 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 161 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 162 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 163 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 164 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 165 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 166 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 167 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 168 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 169 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 170 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 171 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 172 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 173 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 174 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 175 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 176 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 177 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 178 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 179 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 180 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 181 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 182 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 183 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 184 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 185 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 186 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 187 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 188 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 189 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 190 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 191 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 192 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 193 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 194 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 195 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 196 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 197 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 198 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 199 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 200 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 201 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 202 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 203 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 204 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 205 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 206 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 207 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 208 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 209 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 210 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 211 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 212 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 213 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 214 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 215 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 216 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 217 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 218 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 219 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 220 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 221 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 222 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 223 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 224 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 225 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 226 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 227 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 228 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 229 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 230 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 231 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 232 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 233 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 234 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 235 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 236 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 237 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 238 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 239 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 240 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 241 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 242 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 243 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 244 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 245 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 246 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 247 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 248 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 249 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 250 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 251 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 252 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 253 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 254 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 255 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 256 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 257 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 258 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 259 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 260 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 261 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 262 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 263 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 264 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 265 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 266 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 267 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 268 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 269 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 270 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 271 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 272 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 273 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 274 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 275 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 276 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 277 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 278 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 279 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 280 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 281 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 282 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 283 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 284 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 285 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 286 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 287 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 288 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 289 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 290 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 291 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 292 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 293 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 294 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 295 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 296 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 297 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 298 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 299 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 300 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 301 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 302 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 303 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 304 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 305 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 306 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 307 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 308 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 309 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 310 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 311 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 312 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 313 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 314 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 315 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 316 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 317 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 318 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 319 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 320 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 321 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 322 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 323 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 324 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 325 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 326 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 327 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 328 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 329 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 330 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 331 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 332 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 333 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 334 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 335 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 336 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 337 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 338 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 339 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 340 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 341 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 342 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 343 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 344 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 345 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 346 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 347 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 348 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 349 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 350 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 351 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 352 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 353 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 354 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 355 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 356 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 357 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 358 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 359 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 360 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 361 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 362 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 363 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 364 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 365 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 366 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 367 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 368 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 369 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 370 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 371 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 372 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 373 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 374 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 375 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 376 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 377 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 378 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 379 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 380 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 381 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 382 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 383 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 384 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 385 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 386 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 387 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 388 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 389 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 390 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 391 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 392 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 393 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 394 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 395 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 396 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 397 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 398 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 399 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 400 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 401 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 402 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 403 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 404 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 405 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 406 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 407 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 408 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 409 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 410 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 411 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 412 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 413 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 414 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 415 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 416 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 417 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 418 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 419 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 420 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 421 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 422 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 423 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 424 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 425 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 426 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 427 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 428 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 429 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 430 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 431 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 432 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 433 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 434 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 435 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 436 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 437 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 438 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 439 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 440 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 441 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 442 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 443 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 444 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 445 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 446 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 447 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 448 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 449 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 450 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 451 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 452 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 453 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 454 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 455 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 456 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 457 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 458 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 459 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 460 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 461 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 462 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 463 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 464 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 465 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 466 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 467 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 468 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 469 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 470 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 471 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 472 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 473 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 474 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 475 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 476 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 477 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 478 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 479 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 480 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 481 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 482 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 483 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 484 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 485 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 486 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 487 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 488 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 489 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 490 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 491 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 492 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 493 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 494 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 495 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 496 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 497 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 498 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 499 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 500 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 501 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 502 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 503 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 504 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 505 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 506 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 507 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 508 nsew default input
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 509 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 510 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 511 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 512 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 513 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 514 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 515 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 516 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 517 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 518 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 519 nsew default tristate
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 520 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 521 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 522 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 523 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 524 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 525 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 526 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 527 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 528 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 529 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 530 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 531 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 532 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 533 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 534 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 535 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 536 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 537 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 538 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 539 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 540 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 541 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 542 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 543 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 544 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 545 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 546 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 547 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 548 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 549 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 550 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 551 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 552 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 553 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 554 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 555 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 556 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 557 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 558 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 559 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 560 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 561 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 562 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 563 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 564 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 565 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 566 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 567 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 568 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 569 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 570 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 571 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 572 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 573 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 574 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 575 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 576 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 577 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 578 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 579 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 580 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 581 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 582 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 583 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 584 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 585 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 586 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 587 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 588 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 589 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 590 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 591 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 592 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 593 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 594 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 595 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 596 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 597 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 598 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 599 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 600 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 601 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 602 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 603 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 604 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 605 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 606 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 607 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 608 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 609 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 610 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 611 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 612 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 613 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 614 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 615 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 616 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 617 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 618 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 619 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 620 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 621 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 622 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 623 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 624 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 625 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 626 nsew default input
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 627 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 628 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 629 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 630 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 631 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 632 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 633 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 634 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 635 nsew default tristate
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1
port 637 nsew default input
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2
port 638 nsew default input
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2
port 639 nsew default input
rlabel metal5 s -5756 -4684 589680 -4084 8 vdda1
port 640 nsew default input
rlabel metal5 s -6696 -5624 590620 -5024 8 vssa1
port 641 nsew default input
rlabel metal5 s -7636 -6564 591560 -5964 8 vdda2
port 642 nsew default input
rlabel metal5 s -8576 -7504 592500 -6904 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO decred_controller
  CLASS BLOCK ;
  FOREIGN decred_controller ;
  ORIGIN 0.000 0.000 ;
  SIZE 205.000 BY 205.000 ;
  PIN CLK_LED
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 201.000 16.930 205.000 ;
    END
  END CLK_LED
  PIN DATA_AVAILABLE[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 201.000 112.610 205.000 ;
    END
  END DATA_AVAILABLE[0]
  PIN DATA_AVAILABLE[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 201.000 91.450 205.000 ;
    END
  END DATA_AVAILABLE[1]
  PIN DATA_AVAILABLE[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END DATA_AVAILABLE[2]
  PIN DATA_AVAILABLE[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 201.000 176.090 205.000 ;
    END
  END DATA_AVAILABLE[3]
  PIN DATA_FROM_HASH[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END DATA_FROM_HASH[0]
  PIN DATA_FROM_HASH[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END DATA_FROM_HASH[1]
  PIN DATA_FROM_HASH[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 201.000 154.930 205.000 ;
    END
  END DATA_FROM_HASH[2]
  PIN DATA_FROM_HASH[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 201.000 27.970 205.000 ;
    END
  END DATA_FROM_HASH[3]
  PIN DATA_FROM_HASH[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END DATA_FROM_HASH[4]
  PIN DATA_FROM_HASH[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.000 51.720 205.000 52.320 ;
    END
  END DATA_FROM_HASH[5]
  PIN DATA_FROM_HASH[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 201.000 80.410 205.000 ;
    END
  END DATA_FROM_HASH[6]
  PIN DATA_FROM_HASH[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END DATA_FROM_HASH[7]
  PIN DATA_TO_HASH[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END DATA_TO_HASH[0]
  PIN DATA_TO_HASH[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 201.000 186.210 205.000 ;
    END
  END DATA_TO_HASH[1]
  PIN DATA_TO_HASH[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END DATA_TO_HASH[2]
  PIN DATA_TO_HASH[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 0.000 182.530 4.000 ;
    END
  END DATA_TO_HASH[3]
  PIN DATA_TO_HASH[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 201.000 38.090 205.000 ;
    END
  END DATA_TO_HASH[4]
  PIN DATA_TO_HASH[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.000 5.480 205.000 6.080 ;
    END
  END DATA_TO_HASH[5]
  PIN DATA_TO_HASH[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.000 99.320 205.000 99.920 ;
    END
  END DATA_TO_HASH[6]
  PIN DATA_TO_HASH[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 0.000 171.490 4.000 ;
    END
  END DATA_TO_HASH[7]
  PIN EXT_RESET_N_fromHost
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 201.000 122.730 205.000 ;
    END
  END EXT_RESET_N_fromHost
  PIN EXT_RESET_N_toClient
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END EXT_RESET_N_toClient
  PIN HASH_ADDR[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END HASH_ADDR[0]
  PIN HASH_ADDR[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 201.000 165.050 205.000 ;
    END
  END HASH_ADDR[1]
  PIN HASH_ADDR[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END HASH_ADDR[2]
  PIN HASH_ADDR[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 201.000 143.890 205.000 ;
    END
  END HASH_ADDR[3]
  PIN HASH_ADDR[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END HASH_ADDR[4]
  PIN HASH_ADDR[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END HASH_ADDR[5]
  PIN HASH_EN
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 201.000 70.290 205.000 ;
    END
  END HASH_EN
  PIN HASH_LED
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END HASH_LED
  PIN ID_fromClient
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.000 68.040 205.000 68.640 ;
    END
  END ID_fromClient
  PIN ID_toHost
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END ID_toHost
  PIN IRQ_OUT_fromClient
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.000 114.280 205.000 114.880 ;
    END
  END IRQ_OUT_fromClient
  PIN IRQ_OUT_toHost
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END IRQ_OUT_toHost
  PIN M1_CLK_IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END M1_CLK_IN
  PIN M1_CLK_SELECT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 0.000 34.410 4.000 ;
    END
  END M1_CLK_SELECT
  PIN MACRO_RD_SELECT[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.930 0.000 140.210 4.000 ;
    END
  END MACRO_RD_SELECT[0]
  PIN MACRO_RD_SELECT[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 0.000 108.010 4.000 ;
    END
  END MACRO_RD_SELECT[1]
  PIN MACRO_RD_SELECT[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 4.000 ;
    END
  END MACRO_RD_SELECT[2]
  PIN MACRO_RD_SELECT[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END MACRO_RD_SELECT[3]
  PIN MACRO_WR_SELECT[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 201.000 49.130 205.000 ;
    END
  END MACRO_WR_SELECT[0]
  PIN MACRO_WR_SELECT[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END MACRO_WR_SELECT[1]
  PIN MACRO_WR_SELECT[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 201.000 197.250 205.000 ;
    END
  END MACRO_WR_SELECT[2]
  PIN MACRO_WR_SELECT[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.000 36.760 205.000 37.360 ;
    END
  END MACRO_WR_SELECT[3]
  PIN MISO_fromClient
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 201.000 6.810 205.000 ;
    END
  END MISO_fromClient
  PIN MISO_toHost
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 201.000 133.770 205.000 ;
    END
  END MISO_toHost
  PIN MOSI_fromHost
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.000 193.160 205.000 193.760 ;
    END
  END MOSI_fromHost
  PIN MOSI_toClient
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.000 83.000 205.000 83.600 ;
    END
  END MOSI_toClient
  PIN PLL_INPUT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.000 20.440 205.000 21.040 ;
    END
  END PLL_INPUT
  PIN S1_CLK_IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END S1_CLK_IN
  PIN S1_CLK_SELECT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.000 176.840 205.000 177.440 ;
    END
  END S1_CLK_SELECT
  PIN SCLK_fromHost
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.000 161.880 205.000 162.480 ;
    END
  END SCLK_fromHost
  PIN SCLK_toClient
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END SCLK_toClient
  PIN SCSN_fromHost
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 201.000 101.570 205.000 ;
    END
  END SCSN_fromHost
  PIN SCSN_toClient
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.000 145.560 205.000 146.160 ;
    END
  END SCSN_toClient
  PIN THREAD_COUNT[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END THREAD_COUNT[0]
  PIN THREAD_COUNT[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.000 130.600 205.000 131.200 ;
    END
  END THREAD_COUNT[1]
  PIN THREAD_COUNT[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END THREAD_COUNT[2]
  PIN THREAD_COUNT[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 201.000 59.250 205.000 ;
    END
  END THREAD_COUNT[3]
  PIN m1_clk_local
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END m1_clk_local
  PIN one
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END one
  PIN zero
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END zero
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 193.360 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 193.360 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 193.360 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 177.940 10.880 179.540 193.120 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.880 25.940 193.120 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 101.140 10.880 102.740 193.120 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 181.240 10.880 182.840 193.120 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 27.640 10.880 29.240 193.120 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 104.440 10.880 106.040 193.120 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 184.540 10.880 186.140 193.120 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 30.940 10.880 32.540 193.120 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 107.740 10.880 109.340 193.120 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 199.180 193.205 ;
      LAYER met1 ;
        RECT 2.830 8.880 199.180 193.360 ;
      LAYER met2 ;
        RECT 2.860 200.720 6.250 201.000 ;
        RECT 7.090 200.720 16.370 201.000 ;
        RECT 17.210 200.720 27.410 201.000 ;
        RECT 28.250 200.720 37.530 201.000 ;
        RECT 38.370 200.720 48.570 201.000 ;
        RECT 49.410 200.720 58.690 201.000 ;
        RECT 59.530 200.720 69.730 201.000 ;
        RECT 70.570 200.720 79.850 201.000 ;
        RECT 80.690 200.720 90.890 201.000 ;
        RECT 91.730 200.720 101.010 201.000 ;
        RECT 101.850 200.720 112.050 201.000 ;
        RECT 112.890 200.720 122.170 201.000 ;
        RECT 123.010 200.720 133.210 201.000 ;
        RECT 134.050 200.720 143.330 201.000 ;
        RECT 144.170 200.720 154.370 201.000 ;
        RECT 155.210 200.720 164.490 201.000 ;
        RECT 165.330 200.720 175.530 201.000 ;
        RECT 176.370 200.720 185.650 201.000 ;
        RECT 186.490 200.720 196.690 201.000 ;
        RECT 2.860 4.280 197.240 200.720 ;
        RECT 3.410 4.000 12.690 4.280 ;
        RECT 13.530 4.000 22.810 4.280 ;
        RECT 23.650 4.000 33.850 4.280 ;
        RECT 34.690 4.000 43.970 4.280 ;
        RECT 44.810 4.000 55.010 4.280 ;
        RECT 55.850 4.000 65.130 4.280 ;
        RECT 65.970 4.000 76.170 4.280 ;
        RECT 77.010 4.000 86.290 4.280 ;
        RECT 87.130 4.000 97.330 4.280 ;
        RECT 98.170 4.000 107.450 4.280 ;
        RECT 108.290 4.000 118.490 4.280 ;
        RECT 119.330 4.000 128.610 4.280 ;
        RECT 129.450 4.000 139.650 4.280 ;
        RECT 140.490 4.000 149.770 4.280 ;
        RECT 150.610 4.000 160.810 4.280 ;
        RECT 161.650 4.000 170.930 4.280 ;
        RECT 171.770 4.000 181.970 4.280 ;
        RECT 182.810 4.000 192.090 4.280 ;
        RECT 192.930 4.000 197.240 4.280 ;
      LAYER met3 ;
        RECT 4.000 192.760 200.600 193.625 ;
        RECT 4.000 191.440 201.000 192.760 ;
        RECT 4.400 190.040 201.000 191.440 ;
        RECT 4.000 177.840 201.000 190.040 ;
        RECT 4.000 176.480 200.600 177.840 ;
        RECT 4.400 176.440 200.600 176.480 ;
        RECT 4.400 175.080 201.000 176.440 ;
        RECT 4.000 162.880 201.000 175.080 ;
        RECT 4.000 161.480 200.600 162.880 ;
        RECT 4.000 160.160 201.000 161.480 ;
        RECT 4.400 158.760 201.000 160.160 ;
        RECT 4.000 146.560 201.000 158.760 ;
        RECT 4.000 145.200 200.600 146.560 ;
        RECT 4.400 145.160 200.600 145.200 ;
        RECT 4.400 143.800 201.000 145.160 ;
        RECT 4.000 131.600 201.000 143.800 ;
        RECT 4.000 130.200 200.600 131.600 ;
        RECT 4.000 128.880 201.000 130.200 ;
        RECT 4.400 127.480 201.000 128.880 ;
        RECT 4.000 115.280 201.000 127.480 ;
        RECT 4.000 113.920 200.600 115.280 ;
        RECT 4.400 113.880 200.600 113.920 ;
        RECT 4.400 112.520 201.000 113.880 ;
        RECT 4.000 100.320 201.000 112.520 ;
        RECT 4.000 98.920 200.600 100.320 ;
        RECT 4.000 97.600 201.000 98.920 ;
        RECT 4.400 96.200 201.000 97.600 ;
        RECT 4.000 84.000 201.000 96.200 ;
        RECT 4.000 82.640 200.600 84.000 ;
        RECT 4.400 82.600 200.600 82.640 ;
        RECT 4.400 81.240 201.000 82.600 ;
        RECT 4.000 69.040 201.000 81.240 ;
        RECT 4.000 67.640 200.600 69.040 ;
        RECT 4.000 66.320 201.000 67.640 ;
        RECT 4.400 64.920 201.000 66.320 ;
        RECT 4.000 52.720 201.000 64.920 ;
        RECT 4.000 51.360 200.600 52.720 ;
        RECT 4.400 51.320 200.600 51.360 ;
        RECT 4.400 49.960 201.000 51.320 ;
        RECT 4.000 37.760 201.000 49.960 ;
        RECT 4.000 36.360 200.600 37.760 ;
        RECT 4.000 35.040 201.000 36.360 ;
        RECT 4.400 33.640 201.000 35.040 ;
        RECT 4.000 21.440 201.000 33.640 ;
        RECT 4.000 20.080 200.600 21.440 ;
        RECT 4.400 20.040 200.600 20.080 ;
        RECT 4.400 18.680 201.000 20.040 ;
        RECT 4.000 6.480 201.000 18.680 ;
        RECT 4.000 5.615 200.600 6.480 ;
      LAYER met4 ;
        RECT 94.135 115.775 94.465 144.665 ;
  END
END decred_controller
END LIBRARY


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO decred_controller
  CLASS BLOCK ;
  FOREIGN decred_controller ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 200.000 ;
  PIN CLK_LED
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 16.650 196.000 16.930 200.000 ;
    END
  END CLK_LED
  PIN DATA_AVAILABLE[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 109.570 196.000 109.850 200.000 ;
    END
  END DATA_AVAILABLE[0]
  PIN DATA_AVAILABLE[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 88.410 196.000 88.690 200.000 ;
    END
  END DATA_AVAILABLE[1]
  PIN DATA_AVAILABLE[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END DATA_AVAILABLE[2]
  PIN DATA_AVAILABLE[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 171.210 196.000 171.490 200.000 ;
    END
  END DATA_AVAILABLE[3]
  PIN DATA_FROM_HASH[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 4.000 ;
    END
  END DATA_FROM_HASH[0]
  PIN DATA_FROM_HASH[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END DATA_FROM_HASH[1]
  PIN DATA_FROM_HASH[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 150.050 196.000 150.330 200.000 ;
    END
  END DATA_FROM_HASH[2]
  PIN DATA_FROM_HASH[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.770 196.000 27.050 200.000 ;
    END
  END DATA_FROM_HASH[3]
  PIN DATA_FROM_HASH[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END DATA_FROM_HASH[4]
  PIN DATA_FROM_HASH[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 50.360 200.000 50.960 ;
    END
  END DATA_FROM_HASH[5]
  PIN DATA_FROM_HASH[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.290 196.000 78.570 200.000 ;
    END
  END DATA_FROM_HASH[6]
  PIN DATA_FROM_HASH[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END DATA_FROM_HASH[7]
  PIN DATA_TO_HASH[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END DATA_TO_HASH[0]
  PIN DATA_TO_HASH[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 181.330 196.000 181.610 200.000 ;
    END
  END DATA_TO_HASH[1]
  PIN DATA_TO_HASH[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END DATA_TO_HASH[2]
  PIN DATA_TO_HASH[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 176.730 0.000 177.010 4.000 ;
    END
  END DATA_TO_HASH[3]
  PIN DATA_TO_HASH[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 36.890 196.000 37.170 200.000 ;
    END
  END DATA_TO_HASH[4]
  PIN DATA_TO_HASH[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 5.480 200.000 6.080 ;
    END
  END DATA_TO_HASH[5]
  PIN DATA_TO_HASH[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 96.600 200.000 97.200 ;
    END
  END DATA_TO_HASH[6]
  PIN DATA_TO_HASH[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 166.610 0.000 166.890 4.000 ;
    END
  END DATA_TO_HASH[7]
  PIN EXT_RESET_N_fromHost
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 119.690 196.000 119.970 200.000 ;
    END
  END EXT_RESET_N_fromHost
  PIN EXT_RESET_N_toClient
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END EXT_RESET_N_toClient
  PIN HASH_ADDR[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 156.490 0.000 156.770 4.000 ;
    END
  END HASH_ADDR[0]
  PIN HASH_ADDR[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 160.170 196.000 160.450 200.000 ;
    END
  END HASH_ADDR[1]
  PIN HASH_ADDR[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END HASH_ADDR[2]
  PIN HASH_ADDR[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 139.930 196.000 140.210 200.000 ;
    END
  END HASH_ADDR[3]
  PIN HASH_ADDR[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END HASH_ADDR[4]
  PIN HASH_ADDR[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END HASH_ADDR[5]
  PIN HASH_EN
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 68.170 196.000 68.450 200.000 ;
    END
  END HASH_EN
  PIN HASH_LED
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END HASH_LED
  PIN ID_fromClient
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 66.680 200.000 67.280 ;
    END
  END ID_fromClient
  PIN ID_toHost
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END ID_toHost
  PIN IRQ_OUT_fromClient
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 111.560 200.000 112.160 ;
    END
  END IRQ_OUT_fromClient
  PIN IRQ_OUT_toHost
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END IRQ_OUT_toHost
  PIN M1_CLK_IN
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END M1_CLK_IN
  PIN M1_CLK_SELECT
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END M1_CLK_SELECT
  PIN MACRO_RD_SELECT[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 136.250 0.000 136.530 4.000 ;
    END
  END MACRO_RD_SELECT[0]
  PIN MACRO_RD_SELECT[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 4.000 ;
    END
  END MACRO_RD_SELECT[1]
  PIN MACRO_RD_SELECT[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END MACRO_RD_SELECT[2]
  PIN MACRO_RD_SELECT[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END MACRO_RD_SELECT[3]
  PIN MACRO_WR_SELECT[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 47.010 196.000 47.290 200.000 ;
    END
  END MACRO_WR_SELECT[0]
  PIN MACRO_WR_SELECT[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END MACRO_WR_SELECT[1]
  PIN MACRO_WR_SELECT[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 191.450 196.000 191.730 200.000 ;
    END
  END MACRO_WR_SELECT[2]
  PIN MACRO_WR_SELECT[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 35.400 200.000 36.000 ;
    END
  END MACRO_WR_SELECT[3]
  PIN MISO_fromClient
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.530 196.000 6.810 200.000 ;
    END
  END MISO_fromClient
  PIN MISO_toHost
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 129.810 196.000 130.090 200.000 ;
    END
  END MISO_toHost
  PIN MOSI_fromHost
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 187.720 200.000 188.320 ;
    END
  END MOSI_fromHost
  PIN MOSI_toClient
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 81.640 200.000 82.240 ;
    END
  END MOSI_toClient
  PIN PLL_INPUT
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 20.440 200.000 21.040 ;
    END
  END PLL_INPUT
  PIN S1_CLK_IN
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END S1_CLK_IN
  PIN S1_CLK_SELECT
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 172.760 200.000 173.360 ;
    END
  END S1_CLK_SELECT
  PIN SCLK_fromHost
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 157.800 200.000 158.400 ;
    END
  END SCLK_fromHost
  PIN SCLK_toClient
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END SCLK_toClient
  PIN SCSN_fromHost
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 98.530 196.000 98.810 200.000 ;
    END
  END SCSN_fromHost
  PIN SCSN_toClient
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 141.480 200.000 142.080 ;
    END
  END SCSN_toClient
  PIN THREAD_COUNT[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END THREAD_COUNT[0]
  PIN THREAD_COUNT[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 126.520 200.000 127.120 ;
    END
  END THREAD_COUNT[1]
  PIN THREAD_COUNT[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END THREAD_COUNT[2]
  PIN THREAD_COUNT[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.050 196.000 58.330 200.000 ;
    END
  END THREAD_COUNT[3]
  PIN m1_clk_local
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END m1_clk_local
  PIN one
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 146.370 0.000 146.650 4.000 ;
    END
  END one
  PIN zero
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 4.000 ;
    END
  END zero
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 187.920 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 187.920 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 187.765 ;
      LAYER met1 ;
        RECT 5.520 9.560 194.120 195.800 ;
      LAYER met2 ;
        RECT 2.850 195.720 6.250 196.000 ;
        RECT 7.090 195.720 16.370 196.000 ;
        RECT 17.210 195.720 26.490 196.000 ;
        RECT 27.330 195.720 36.610 196.000 ;
        RECT 37.450 195.720 46.730 196.000 ;
        RECT 47.570 195.720 57.770 196.000 ;
        RECT 58.610 195.720 67.890 196.000 ;
        RECT 68.730 195.720 78.010 196.000 ;
        RECT 78.850 195.720 88.130 196.000 ;
        RECT 88.970 195.720 98.250 196.000 ;
        RECT 99.090 195.720 109.290 196.000 ;
        RECT 110.130 195.720 119.410 196.000 ;
        RECT 120.250 195.720 129.530 196.000 ;
        RECT 130.370 195.720 139.650 196.000 ;
        RECT 140.490 195.720 149.770 196.000 ;
        RECT 150.610 195.720 159.890 196.000 ;
        RECT 160.730 195.720 170.930 196.000 ;
        RECT 171.770 195.720 181.050 196.000 ;
        RECT 181.890 195.720 191.170 196.000 ;
        RECT 2.850 4.280 191.720 195.720 ;
        RECT 3.410 4.000 12.690 4.280 ;
        RECT 13.530 4.000 22.810 4.280 ;
        RECT 23.650 4.000 32.930 4.280 ;
        RECT 33.770 4.000 43.050 4.280 ;
        RECT 43.890 4.000 53.170 4.280 ;
        RECT 54.010 4.000 64.210 4.280 ;
        RECT 65.050 4.000 74.330 4.280 ;
        RECT 75.170 4.000 84.450 4.280 ;
        RECT 85.290 4.000 94.570 4.280 ;
        RECT 95.410 4.000 104.690 4.280 ;
        RECT 105.530 4.000 114.810 4.280 ;
        RECT 115.650 4.000 125.850 4.280 ;
        RECT 126.690 4.000 135.970 4.280 ;
        RECT 136.810 4.000 146.090 4.280 ;
        RECT 146.930 4.000 156.210 4.280 ;
        RECT 157.050 4.000 166.330 4.280 ;
        RECT 167.170 4.000 176.450 4.280 ;
        RECT 177.290 4.000 187.490 4.280 ;
        RECT 188.330 4.000 191.720 4.280 ;
      LAYER met3 ;
        RECT 2.825 187.360 195.600 188.185 ;
        RECT 4.400 187.320 195.600 187.360 ;
        RECT 4.400 185.960 196.000 187.320 ;
        RECT 2.825 173.760 196.000 185.960 ;
        RECT 2.825 172.360 195.600 173.760 ;
        RECT 2.825 171.040 196.000 172.360 ;
        RECT 4.400 169.640 196.000 171.040 ;
        RECT 2.825 158.800 196.000 169.640 ;
        RECT 2.825 157.400 195.600 158.800 ;
        RECT 2.825 156.080 196.000 157.400 ;
        RECT 4.400 154.680 196.000 156.080 ;
        RECT 2.825 142.480 196.000 154.680 ;
        RECT 2.825 141.120 195.600 142.480 ;
        RECT 4.400 141.080 195.600 141.120 ;
        RECT 4.400 139.720 196.000 141.080 ;
        RECT 2.825 127.520 196.000 139.720 ;
        RECT 2.825 126.160 195.600 127.520 ;
        RECT 4.400 126.120 195.600 126.160 ;
        RECT 4.400 124.760 196.000 126.120 ;
        RECT 2.825 112.560 196.000 124.760 ;
        RECT 2.825 111.200 195.600 112.560 ;
        RECT 4.400 111.160 195.600 111.200 ;
        RECT 4.400 109.800 196.000 111.160 ;
        RECT 2.825 97.600 196.000 109.800 ;
        RECT 2.825 96.240 195.600 97.600 ;
        RECT 4.400 96.200 195.600 96.240 ;
        RECT 4.400 94.840 196.000 96.200 ;
        RECT 2.825 82.640 196.000 94.840 ;
        RECT 2.825 81.240 195.600 82.640 ;
        RECT 2.825 79.920 196.000 81.240 ;
        RECT 4.400 78.520 196.000 79.920 ;
        RECT 2.825 67.680 196.000 78.520 ;
        RECT 2.825 66.280 195.600 67.680 ;
        RECT 2.825 64.960 196.000 66.280 ;
        RECT 4.400 63.560 196.000 64.960 ;
        RECT 2.825 51.360 196.000 63.560 ;
        RECT 2.825 50.000 195.600 51.360 ;
        RECT 4.400 49.960 195.600 50.000 ;
        RECT 4.400 48.600 196.000 49.960 ;
        RECT 2.825 36.400 196.000 48.600 ;
        RECT 2.825 35.040 195.600 36.400 ;
        RECT 4.400 35.000 195.600 35.040 ;
        RECT 4.400 33.640 196.000 35.000 ;
        RECT 2.825 21.440 196.000 33.640 ;
        RECT 2.825 20.080 195.600 21.440 ;
        RECT 4.400 20.040 195.600 20.080 ;
        RECT 4.400 18.680 196.000 20.040 ;
        RECT 2.825 6.480 196.000 18.680 ;
        RECT 2.825 5.615 195.600 6.480 ;
      LAYER met4 ;
        RECT 121.735 10.640 176.240 187.920 ;
  END
END decred_controller
END LIBRARY


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO decred_hash_macro
  CLASS BLOCK ;
  FOREIGN decred_hash_macro ;
  ORIGIN 0.000 0.000 ;
  SIZE 1220.000 BY 1020.000 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.250 1016.000 665.530 1020.000 ;
    END
  END CLK
  PIN DATA_AVAILABLE
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.010 0.000 737.290 4.000 ;
    END
  END DATA_AVAILABLE
  PIN DATA_FROM_HASH[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 0.000 125.490 4.000 ;
    END
  END DATA_FROM_HASH[0]
  PIN DATA_FROM_HASH[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END DATA_FROM_HASH[1]
  PIN DATA_FROM_HASH[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 910.890 1016.000 911.170 1020.000 ;
    END
  END DATA_FROM_HASH[2]
  PIN DATA_FROM_HASH[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1105.010 0.000 1105.290 4.000 ;
    END
  END DATA_FROM_HASH[3]
  PIN DATA_FROM_HASH[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1216.000 199.960 1220.000 200.560 ;
    END
  END DATA_FROM_HASH[4]
  PIN DATA_FROM_HASH[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.930 0.000 370.210 4.000 ;
    END
  END DATA_FROM_HASH[5]
  PIN DATA_FROM_HASH[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 1016.000 176.090 1020.000 ;
    END
  END DATA_FROM_HASH[6]
  PIN DATA_FROM_HASH[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 727.640 4.000 728.240 ;
    END
  END DATA_FROM_HASH[7]
  PIN DATA_TO_HASH[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.530 1016.000 420.810 1020.000 ;
    END
  END DATA_TO_HASH[0]
  PIN DATA_TO_HASH[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.880 4.000 366.480 ;
    END
  END DATA_TO_HASH[1]
  PIN DATA_TO_HASH[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1216.000 380.840 1220.000 381.440 ;
    END
  END DATA_TO_HASH[2]
  PIN DATA_TO_HASH[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1216.000 19.080 1220.000 19.680 ;
    END
  END DATA_TO_HASH[3]
  PIN DATA_TO_HASH[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 908.520 4.000 909.120 ;
    END
  END DATA_TO_HASH[4]
  PIN DATA_TO_HASH[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.570 0.000 247.850 4.000 ;
    END
  END DATA_TO_HASH[5]
  PIN DATA_TO_HASH[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.250 1016.000 1033.530 1020.000 ;
    END
  END DATA_TO_HASH[6]
  PIN DATA_TO_HASH[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 1016.000 298.450 1020.000 ;
    END
  END DATA_TO_HASH[7]
  PIN HASH_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.610 1016.000 787.890 1020.000 ;
    END
  END HASH_ADDR[0]
  PIN HASH_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 1016.000 52.810 1020.000 ;
    END
  END HASH_ADDR[1]
  PIN HASH_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1155.610 1016.000 1155.890 1020.000 ;
    END
  END HASH_ADDR[2]
  PIN HASH_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.650 0.000 982.930 4.000 ;
    END
  END HASH_ADDR[3]
  PIN HASH_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END HASH_ADDR[4]
  PIN HASH_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1216.000 924.840 1220.000 925.440 ;
    END
  END HASH_ADDR[5]
  PIN HASH_EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.290 0.000 492.570 4.000 ;
    END
  END HASH_EN
  PIN MACRO_RD_SELECT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.650 0.000 614.930 4.000 ;
    END
  END MACRO_RD_SELECT
  PIN MACRO_WR_SELECT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1216.000 563.080 1220.000 563.680 ;
    END
  END MACRO_WR_SELECT
  PIN THREAD_COUNT[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1216.000 743.960 1220.000 744.560 ;
    END
  END THREAD_COUNT[0]
  PIN THREAD_COUNT[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 546.760 4.000 547.360 ;
    END
  END THREAD_COUNT[1]
  PIN THREAD_COUNT[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.890 1016.000 543.170 1020.000 ;
    END
  END THREAD_COUNT[2]
  PIN THREAD_COUNT[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.290 0.000 860.570 4.000 ;
    END
  END THREAD_COUNT[3]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1009.360 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1009.360 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1009.360 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1009.360 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1009.360 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1009.360 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1009.360 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1009.360 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1009.360 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1009.360 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1009.360 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1009.360 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1009.360 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1009.360 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1009.360 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1009.360 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1099.540 10.880 1101.140 1009.120 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 945.940 10.880 947.540 1009.120 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 792.340 10.880 793.940 1009.120 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 638.740 10.880 640.340 1009.120 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 485.140 10.880 486.740 1009.120 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 331.540 10.880 333.140 1009.120 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 177.940 10.880 179.540 1009.120 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.880 25.940 1009.120 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1176.340 10.880 1177.940 1009.120 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1022.740 10.880 1024.340 1009.120 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 869.140 10.880 870.740 1009.120 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 715.540 10.880 717.140 1009.120 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 561.940 10.880 563.540 1009.120 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 408.340 10.880 409.940 1009.120 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 254.740 10.880 256.340 1009.120 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 101.140 10.880 102.740 1009.120 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1102.840 10.880 1104.440 1009.120 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 949.240 10.880 950.840 1009.120 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 795.640 10.880 797.240 1009.120 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 642.040 10.880 643.640 1009.120 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 488.440 10.880 490.040 1009.120 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 334.840 10.880 336.440 1009.120 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 181.240 10.880 182.840 1009.120 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 27.640 10.880 29.240 1009.120 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1179.640 10.880 1181.240 1009.120 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1026.040 10.880 1027.640 1009.120 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 872.440 10.880 874.040 1009.120 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 718.840 10.880 720.440 1009.120 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 565.240 10.880 566.840 1009.120 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 411.640 10.880 413.240 1009.120 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 258.040 10.880 259.640 1009.120 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 104.440 10.880 106.040 1009.120 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1106.140 10.880 1107.740 1009.120 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 952.540 10.880 954.140 1009.120 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 798.940 10.880 800.540 1009.120 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 645.340 10.880 646.940 1009.120 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 491.740 10.880 493.340 1009.120 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 338.140 10.880 339.740 1009.120 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 184.540 10.880 186.140 1009.120 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 30.940 10.880 32.540 1009.120 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1182.940 10.880 1184.540 1009.120 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1029.340 10.880 1030.940 1009.120 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 875.740 10.880 877.340 1009.120 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 722.140 10.880 723.740 1009.120 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 568.540 10.880 570.140 1009.120 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 414.940 10.880 416.540 1009.120 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 261.340 10.880 262.940 1009.120 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 107.740 10.880 109.340 1009.120 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1214.400 1009.205 ;
      LAYER met1 ;
        RECT 1.910 8.880 1214.400 1009.360 ;
      LAYER met2 ;
        RECT 1.930 1015.720 52.250 1016.000 ;
        RECT 53.090 1015.720 175.530 1016.000 ;
        RECT 176.370 1015.720 297.890 1016.000 ;
        RECT 298.730 1015.720 420.250 1016.000 ;
        RECT 421.090 1015.720 542.610 1016.000 ;
        RECT 543.450 1015.720 664.970 1016.000 ;
        RECT 665.810 1015.720 787.330 1016.000 ;
        RECT 788.170 1015.720 910.610 1016.000 ;
        RECT 911.450 1015.720 1032.970 1016.000 ;
        RECT 1033.810 1015.720 1155.330 1016.000 ;
        RECT 1156.170 1015.720 1210.630 1016.000 ;
        RECT 1.930 4.280 1210.630 1015.720 ;
        RECT 1.930 4.000 2.570 4.280 ;
        RECT 3.410 4.000 124.930 4.280 ;
        RECT 125.770 4.000 247.290 4.280 ;
        RECT 248.130 4.000 369.650 4.280 ;
        RECT 370.490 4.000 492.010 4.280 ;
        RECT 492.850 4.000 614.370 4.280 ;
        RECT 615.210 4.000 736.730 4.280 ;
        RECT 737.570 4.000 860.010 4.280 ;
        RECT 860.850 4.000 982.370 4.280 ;
        RECT 983.210 4.000 1104.730 4.280 ;
        RECT 1105.570 4.000 1210.630 4.280 ;
      LAYER met3 ;
        RECT 1.905 925.840 1216.000 1009.285 ;
        RECT 1.905 924.440 1215.600 925.840 ;
        RECT 1.905 909.520 1216.000 924.440 ;
        RECT 4.400 908.120 1216.000 909.520 ;
        RECT 1.905 744.960 1216.000 908.120 ;
        RECT 1.905 743.560 1215.600 744.960 ;
        RECT 1.905 728.640 1216.000 743.560 ;
        RECT 4.400 727.240 1216.000 728.640 ;
        RECT 1.905 564.080 1216.000 727.240 ;
        RECT 1.905 562.680 1215.600 564.080 ;
        RECT 1.905 547.760 1216.000 562.680 ;
        RECT 4.400 546.360 1216.000 547.760 ;
        RECT 1.905 381.840 1216.000 546.360 ;
        RECT 1.905 380.440 1215.600 381.840 ;
        RECT 1.905 366.880 1216.000 380.440 ;
        RECT 4.400 365.480 1216.000 366.880 ;
        RECT 1.905 200.960 1216.000 365.480 ;
        RECT 1.905 199.560 1215.600 200.960 ;
        RECT 1.905 186.000 1216.000 199.560 ;
        RECT 4.400 184.600 1216.000 186.000 ;
        RECT 1.905 20.080 1216.000 184.600 ;
        RECT 1.905 18.680 1215.600 20.080 ;
        RECT 1.905 10.715 1216.000 18.680 ;
      LAYER met4 ;
        RECT 3.055 16.495 20.640 1004.865 ;
        RECT 23.040 16.495 23.940 1004.865 ;
        RECT 26.340 16.495 27.240 1004.865 ;
        RECT 29.640 16.495 30.540 1004.865 ;
        RECT 32.940 16.495 97.440 1004.865 ;
        RECT 99.840 16.495 100.740 1004.865 ;
        RECT 103.140 16.495 104.040 1004.865 ;
        RECT 106.440 16.495 107.340 1004.865 ;
        RECT 109.740 16.495 174.240 1004.865 ;
        RECT 176.640 16.495 177.540 1004.865 ;
        RECT 179.940 16.495 180.840 1004.865 ;
        RECT 183.240 16.495 184.140 1004.865 ;
        RECT 186.540 16.495 251.040 1004.865 ;
        RECT 253.440 16.495 254.340 1004.865 ;
        RECT 256.740 16.495 257.640 1004.865 ;
        RECT 260.040 16.495 260.940 1004.865 ;
        RECT 263.340 16.495 327.840 1004.865 ;
        RECT 330.240 16.495 331.140 1004.865 ;
        RECT 333.540 16.495 334.440 1004.865 ;
        RECT 336.840 16.495 337.740 1004.865 ;
        RECT 340.140 16.495 404.640 1004.865 ;
        RECT 407.040 16.495 407.940 1004.865 ;
        RECT 410.340 16.495 411.240 1004.865 ;
        RECT 413.640 16.495 414.540 1004.865 ;
        RECT 416.940 16.495 481.440 1004.865 ;
        RECT 483.840 16.495 484.740 1004.865 ;
        RECT 487.140 16.495 488.040 1004.865 ;
        RECT 490.440 16.495 491.340 1004.865 ;
        RECT 493.740 16.495 558.240 1004.865 ;
        RECT 560.640 16.495 561.540 1004.865 ;
        RECT 563.940 16.495 564.840 1004.865 ;
        RECT 567.240 16.495 568.140 1004.865 ;
        RECT 570.540 16.495 635.040 1004.865 ;
        RECT 637.440 16.495 638.340 1004.865 ;
        RECT 640.740 16.495 641.640 1004.865 ;
        RECT 644.040 16.495 644.940 1004.865 ;
        RECT 647.340 16.495 711.840 1004.865 ;
        RECT 714.240 16.495 715.140 1004.865 ;
        RECT 717.540 16.495 718.440 1004.865 ;
        RECT 720.840 16.495 721.740 1004.865 ;
        RECT 724.140 16.495 788.640 1004.865 ;
        RECT 791.040 16.495 791.940 1004.865 ;
        RECT 794.340 16.495 795.240 1004.865 ;
        RECT 797.640 16.495 798.540 1004.865 ;
        RECT 800.940 16.495 865.440 1004.865 ;
        RECT 867.840 16.495 868.740 1004.865 ;
        RECT 871.140 16.495 872.040 1004.865 ;
        RECT 874.440 16.495 875.340 1004.865 ;
        RECT 877.740 16.495 942.240 1004.865 ;
        RECT 944.640 16.495 945.540 1004.865 ;
        RECT 947.940 16.495 948.840 1004.865 ;
        RECT 951.240 16.495 952.140 1004.865 ;
        RECT 954.540 16.495 1019.040 1004.865 ;
        RECT 1021.440 16.495 1022.340 1004.865 ;
        RECT 1024.740 16.495 1025.640 1004.865 ;
        RECT 1028.040 16.495 1028.940 1004.865 ;
        RECT 1031.340 16.495 1095.840 1004.865 ;
        RECT 1098.240 16.495 1099.140 1004.865 ;
        RECT 1101.540 16.495 1102.440 1004.865 ;
        RECT 1104.840 16.495 1105.740 1004.865 ;
        RECT 1108.140 16.495 1172.640 1004.865 ;
        RECT 1175.040 16.495 1175.940 1004.865 ;
        RECT 1178.340 16.495 1179.240 1004.865 ;
        RECT 1181.640 16.495 1182.540 1004.865 ;
        RECT 1184.940 16.495 1196.625 1004.865 ;
      LAYER met5 ;
        RECT 765.100 731.900 808.100 740.300 ;
  END
END decred_hash_macro
END LIBRARY

